magic
tech EFXH018D
magscale 1 2
timestamp 1533305873
<< mimcap >>
rect -38335 6130 -34335 6160
rect -38335 190 -38305 6130
rect -34365 190 -34335 6130
rect -38335 160 -34335 190
rect -33805 6130 -29805 6160
rect -33805 190 -33775 6130
rect -29835 190 -29805 6130
rect -33805 160 -29805 190
rect -29275 6130 -25275 6160
rect -29275 190 -29245 6130
rect -25305 190 -25275 6130
rect -29275 160 -25275 190
rect -24745 6130 -20745 6160
rect -24745 190 -24715 6130
rect -20775 190 -20745 6130
rect -24745 160 -20745 190
rect -20215 6130 -16215 6160
rect -20215 190 -20185 6130
rect -16245 190 -16215 6130
rect -20215 160 -16215 190
rect -15685 6130 -11685 6160
rect -15685 190 -15655 6130
rect -11715 190 -11685 6130
rect -15685 160 -11685 190
rect -11155 6130 -7155 6160
rect -11155 190 -11125 6130
rect -7185 190 -7155 6130
rect -11155 160 -7155 190
rect -6625 6130 -2625 6160
rect -6625 190 -6595 6130
rect -2655 190 -2625 6130
rect -6625 160 -2625 190
rect -2095 6130 1905 6160
rect -2095 190 -2065 6130
rect 1875 190 1905 6130
rect -2095 160 1905 190
rect 2435 6130 6435 6160
rect 2435 190 2465 6130
rect 6405 190 6435 6130
rect 2435 160 6435 190
rect 6965 6130 10965 6160
rect 6965 190 6995 6130
rect 10935 190 10965 6130
rect 6965 160 10965 190
rect 11495 6130 15495 6160
rect 11495 190 11525 6130
rect 15465 190 15495 6130
rect 11495 160 15495 190
rect 16025 6130 20025 6160
rect 16025 190 16055 6130
rect 19995 190 20025 6130
rect 16025 160 20025 190
rect 20555 6130 24555 6160
rect 20555 190 20585 6130
rect 24525 190 24555 6130
rect 20555 160 24555 190
rect 25085 6130 29085 6160
rect 25085 190 25115 6130
rect 29055 190 29085 6130
rect 25085 160 29085 190
rect 29615 6130 33615 6160
rect 29615 190 29645 6130
rect 33585 190 33615 6130
rect 29615 160 33615 190
rect 34145 6130 38145 6160
rect 34145 190 34175 6130
rect 38115 190 38145 6130
rect 34145 160 38145 190
rect -38335 -190 -34335 -160
rect -38335 -6130 -38305 -190
rect -34365 -6130 -34335 -190
rect -38335 -6160 -34335 -6130
rect -33805 -190 -29805 -160
rect -33805 -6130 -33775 -190
rect -29835 -6130 -29805 -190
rect -33805 -6160 -29805 -6130
rect -29275 -190 -25275 -160
rect -29275 -6130 -29245 -190
rect -25305 -6130 -25275 -190
rect -29275 -6160 -25275 -6130
rect -24745 -190 -20745 -160
rect -24745 -6130 -24715 -190
rect -20775 -6130 -20745 -190
rect -24745 -6160 -20745 -6130
rect -20215 -190 -16215 -160
rect -20215 -6130 -20185 -190
rect -16245 -6130 -16215 -190
rect -20215 -6160 -16215 -6130
rect -15685 -190 -11685 -160
rect -15685 -6130 -15655 -190
rect -11715 -6130 -11685 -190
rect -15685 -6160 -11685 -6130
rect -11155 -190 -7155 -160
rect -11155 -6130 -11125 -190
rect -7185 -6130 -7155 -190
rect -11155 -6160 -7155 -6130
rect -6625 -190 -2625 -160
rect -6625 -6130 -6595 -190
rect -2655 -6130 -2625 -190
rect -6625 -6160 -2625 -6130
rect -2095 -190 1905 -160
rect -2095 -6130 -2065 -190
rect 1875 -6130 1905 -190
rect -2095 -6160 1905 -6130
rect 2435 -190 6435 -160
rect 2435 -6130 2465 -190
rect 6405 -6130 6435 -190
rect 2435 -6160 6435 -6130
rect 6965 -190 10965 -160
rect 6965 -6130 6995 -190
rect 10935 -6130 10965 -190
rect 6965 -6160 10965 -6130
rect 11495 -190 15495 -160
rect 11495 -6130 11525 -190
rect 15465 -6130 15495 -190
rect 11495 -6160 15495 -6130
rect 16025 -190 20025 -160
rect 16025 -6130 16055 -190
rect 19995 -6130 20025 -190
rect 16025 -6160 20025 -6130
rect 20555 -190 24555 -160
rect 20555 -6130 20585 -190
rect 24525 -6130 24555 -190
rect 20555 -6160 24555 -6130
rect 25085 -190 29085 -160
rect 25085 -6130 25115 -190
rect 29055 -6130 29085 -190
rect 25085 -6160 29085 -6130
rect 29615 -190 33615 -160
rect 29615 -6130 29645 -190
rect 33585 -6130 33615 -190
rect 29615 -6160 33615 -6130
rect 34145 -190 38145 -160
rect 34145 -6130 34175 -190
rect 38115 -6130 38145 -190
rect 34145 -6160 38145 -6130
<< mimcapcontact >>
rect -38305 190 -34365 6130
rect -33775 190 -29835 6130
rect -29245 190 -25305 6130
rect -24715 190 -20775 6130
rect -20185 190 -16245 6130
rect -15655 190 -11715 6130
rect -11125 190 -7185 6130
rect -6595 190 -2655 6130
rect -2065 190 1875 6130
rect 2465 190 6405 6130
rect 6995 190 10935 6130
rect 11525 190 15465 6130
rect 16055 190 19995 6130
rect 20585 190 24525 6130
rect 25115 190 29055 6130
rect 29645 190 33585 6130
rect 34175 190 38115 6130
rect -38305 -6130 -34365 -190
rect -33775 -6130 -29835 -190
rect -29245 -6130 -25305 -190
rect -24715 -6130 -20775 -190
rect -20185 -6130 -16245 -190
rect -15655 -6130 -11715 -190
rect -11125 -6130 -7185 -190
rect -6595 -6130 -2655 -190
rect -2065 -6130 1875 -190
rect 2465 -6130 6405 -190
rect 6995 -6130 10935 -190
rect 11525 -6130 15465 -190
rect 16055 -6130 19995 -190
rect 20585 -6130 24525 -190
rect 25115 -6130 29055 -190
rect 29645 -6130 33585 -190
rect 34175 -6130 38115 -190
<< metal4 >>
rect -38435 6232 -34045 6260
rect -38435 6160 -34165 6232
rect -38435 160 -38335 6160
rect -34335 160 -34165 6160
rect -38435 88 -34165 160
rect -34065 88 -34045 6232
rect -38435 60 -34045 88
rect -33905 6232 -29515 6260
rect -33905 6160 -29635 6232
rect -33905 160 -33805 6160
rect -29805 160 -29635 6160
rect -33905 88 -29635 160
rect -29535 88 -29515 6232
rect -33905 60 -29515 88
rect -29375 6232 -24985 6260
rect -29375 6160 -25105 6232
rect -29375 160 -29275 6160
rect -25275 160 -25105 6160
rect -29375 88 -25105 160
rect -25005 88 -24985 6232
rect -29375 60 -24985 88
rect -24845 6232 -20455 6260
rect -24845 6160 -20575 6232
rect -24845 160 -24745 6160
rect -20745 160 -20575 6160
rect -24845 88 -20575 160
rect -20475 88 -20455 6232
rect -24845 60 -20455 88
rect -20315 6232 -15925 6260
rect -20315 6160 -16045 6232
rect -20315 160 -20215 6160
rect -16215 160 -16045 6160
rect -20315 88 -16045 160
rect -15945 88 -15925 6232
rect -20315 60 -15925 88
rect -15785 6232 -11395 6260
rect -15785 6160 -11515 6232
rect -15785 160 -15685 6160
rect -11685 160 -11515 6160
rect -15785 88 -11515 160
rect -11415 88 -11395 6232
rect -15785 60 -11395 88
rect -11255 6232 -6865 6260
rect -11255 6160 -6985 6232
rect -11255 160 -11155 6160
rect -7155 160 -6985 6160
rect -11255 88 -6985 160
rect -6885 88 -6865 6232
rect -11255 60 -6865 88
rect -6725 6232 -2335 6260
rect -6725 6160 -2455 6232
rect -6725 160 -6625 6160
rect -2625 160 -2455 6160
rect -6725 88 -2455 160
rect -2355 88 -2335 6232
rect -6725 60 -2335 88
rect -2195 6232 2195 6260
rect -2195 6160 2075 6232
rect -2195 160 -2095 6160
rect 1905 160 2075 6160
rect -2195 88 2075 160
rect 2175 88 2195 6232
rect -2195 60 2195 88
rect 2335 6232 6725 6260
rect 2335 6160 6605 6232
rect 2335 160 2435 6160
rect 6435 160 6605 6160
rect 2335 88 6605 160
rect 6705 88 6725 6232
rect 2335 60 6725 88
rect 6865 6232 11255 6260
rect 6865 6160 11135 6232
rect 6865 160 6965 6160
rect 10965 160 11135 6160
rect 6865 88 11135 160
rect 11235 88 11255 6232
rect 6865 60 11255 88
rect 11395 6232 15785 6260
rect 11395 6160 15665 6232
rect 11395 160 11495 6160
rect 15495 160 15665 6160
rect 11395 88 15665 160
rect 15765 88 15785 6232
rect 11395 60 15785 88
rect 15925 6232 20315 6260
rect 15925 6160 20195 6232
rect 15925 160 16025 6160
rect 20025 160 20195 6160
rect 15925 88 20195 160
rect 20295 88 20315 6232
rect 15925 60 20315 88
rect 20455 6232 24845 6260
rect 20455 6160 24725 6232
rect 20455 160 20555 6160
rect 24555 160 24725 6160
rect 20455 88 24725 160
rect 24825 88 24845 6232
rect 20455 60 24845 88
rect 24985 6232 29375 6260
rect 24985 6160 29255 6232
rect 24985 160 25085 6160
rect 29085 160 29255 6160
rect 24985 88 29255 160
rect 29355 88 29375 6232
rect 24985 60 29375 88
rect 29515 6232 33905 6260
rect 29515 6160 33785 6232
rect 29515 160 29615 6160
rect 33615 160 33785 6160
rect 29515 88 33785 160
rect 33885 88 33905 6232
rect 29515 60 33905 88
rect 34045 6232 38435 6260
rect 34045 6160 38315 6232
rect 34045 160 34145 6160
rect 38145 160 38315 6160
rect 34045 88 38315 160
rect 38415 88 38435 6232
rect 34045 60 38435 88
rect -38435 -88 -34045 -60
rect -38435 -160 -34165 -88
rect -38435 -6160 -38335 -160
rect -34335 -6160 -34165 -160
rect -38435 -6232 -34165 -6160
rect -34065 -6232 -34045 -88
rect -38435 -6260 -34045 -6232
rect -33905 -88 -29515 -60
rect -33905 -160 -29635 -88
rect -33905 -6160 -33805 -160
rect -29805 -6160 -29635 -160
rect -33905 -6232 -29635 -6160
rect -29535 -6232 -29515 -88
rect -33905 -6260 -29515 -6232
rect -29375 -88 -24985 -60
rect -29375 -160 -25105 -88
rect -29375 -6160 -29275 -160
rect -25275 -6160 -25105 -160
rect -29375 -6232 -25105 -6160
rect -25005 -6232 -24985 -88
rect -29375 -6260 -24985 -6232
rect -24845 -88 -20455 -60
rect -24845 -160 -20575 -88
rect -24845 -6160 -24745 -160
rect -20745 -6160 -20575 -160
rect -24845 -6232 -20575 -6160
rect -20475 -6232 -20455 -88
rect -24845 -6260 -20455 -6232
rect -20315 -88 -15925 -60
rect -20315 -160 -16045 -88
rect -20315 -6160 -20215 -160
rect -16215 -6160 -16045 -160
rect -20315 -6232 -16045 -6160
rect -15945 -6232 -15925 -88
rect -20315 -6260 -15925 -6232
rect -15785 -88 -11395 -60
rect -15785 -160 -11515 -88
rect -15785 -6160 -15685 -160
rect -11685 -6160 -11515 -160
rect -15785 -6232 -11515 -6160
rect -11415 -6232 -11395 -88
rect -15785 -6260 -11395 -6232
rect -11255 -88 -6865 -60
rect -11255 -160 -6985 -88
rect -11255 -6160 -11155 -160
rect -7155 -6160 -6985 -160
rect -11255 -6232 -6985 -6160
rect -6885 -6232 -6865 -88
rect -11255 -6260 -6865 -6232
rect -6725 -88 -2335 -60
rect -6725 -160 -2455 -88
rect -6725 -6160 -6625 -160
rect -2625 -6160 -2455 -160
rect -6725 -6232 -2455 -6160
rect -2355 -6232 -2335 -88
rect -6725 -6260 -2335 -6232
rect -2195 -88 2195 -60
rect -2195 -160 2075 -88
rect -2195 -6160 -2095 -160
rect 1905 -6160 2075 -160
rect -2195 -6232 2075 -6160
rect 2175 -6232 2195 -88
rect -2195 -6260 2195 -6232
rect 2335 -88 6725 -60
rect 2335 -160 6605 -88
rect 2335 -6160 2435 -160
rect 6435 -6160 6605 -160
rect 2335 -6232 6605 -6160
rect 6705 -6232 6725 -88
rect 2335 -6260 6725 -6232
rect 6865 -88 11255 -60
rect 6865 -160 11135 -88
rect 6865 -6160 6965 -160
rect 10965 -6160 11135 -160
rect 6865 -6232 11135 -6160
rect 11235 -6232 11255 -88
rect 6865 -6260 11255 -6232
rect 11395 -88 15785 -60
rect 11395 -160 15665 -88
rect 11395 -6160 11495 -160
rect 15495 -6160 15665 -160
rect 11395 -6232 15665 -6160
rect 15765 -6232 15785 -88
rect 11395 -6260 15785 -6232
rect 15925 -88 20315 -60
rect 15925 -160 20195 -88
rect 15925 -6160 16025 -160
rect 20025 -6160 20195 -160
rect 15925 -6232 20195 -6160
rect 20295 -6232 20315 -88
rect 15925 -6260 20315 -6232
rect 20455 -88 24845 -60
rect 20455 -160 24725 -88
rect 20455 -6160 20555 -160
rect 24555 -6160 24725 -160
rect 20455 -6232 24725 -6160
rect 24825 -6232 24845 -88
rect 20455 -6260 24845 -6232
rect 24985 -88 29375 -60
rect 24985 -160 29255 -88
rect 24985 -6160 25085 -160
rect 29085 -6160 29255 -160
rect 24985 -6232 29255 -6160
rect 29355 -6232 29375 -88
rect 24985 -6260 29375 -6232
rect 29515 -88 33905 -60
rect 29515 -160 33785 -88
rect 29515 -6160 29615 -160
rect 33615 -6160 33785 -160
rect 29515 -6232 33785 -6160
rect 33885 -6232 33905 -88
rect 29515 -6260 33905 -6232
rect 34045 -88 38435 -60
rect 34045 -160 38315 -88
rect 34045 -6160 34145 -160
rect 38145 -6160 38315 -160
rect 34045 -6232 38315 -6160
rect 38415 -6232 38435 -88
rect 34045 -6260 38435 -6232
<< viatp >>
rect -34165 88 -34065 6232
rect -29635 88 -29535 6232
rect -25105 88 -25005 6232
rect -20575 88 -20475 6232
rect -16045 88 -15945 6232
rect -11515 88 -11415 6232
rect -6985 88 -6885 6232
rect -2455 88 -2355 6232
rect 2075 88 2175 6232
rect 6605 88 6705 6232
rect 11135 88 11235 6232
rect 15665 88 15765 6232
rect 20195 88 20295 6232
rect 24725 88 24825 6232
rect 29255 88 29355 6232
rect 33785 88 33885 6232
rect 38315 88 38415 6232
rect -34165 -6232 -34065 -88
rect -29635 -6232 -29535 -88
rect -25105 -6232 -25005 -88
rect -20575 -6232 -20475 -88
rect -16045 -6232 -15945 -88
rect -11515 -6232 -11415 -88
rect -6985 -6232 -6885 -88
rect -2455 -6232 -2355 -88
rect 2075 -6232 2175 -88
rect 6605 -6232 6705 -88
rect 11135 -6232 11235 -88
rect 15665 -6232 15765 -88
rect 20195 -6232 20295 -88
rect 24725 -6232 24825 -88
rect 29255 -6232 29355 -88
rect 33785 -6232 33885 -88
rect 38315 -6232 38415 -88
<< metaltp >>
rect -36405 6130 -36265 6320
rect -34185 6232 -34045 6320
rect -36405 -190 -36265 190
rect -34185 88 -34165 6232
rect -34065 88 -34045 6232
rect -31875 6130 -31735 6320
rect -29655 6232 -29515 6320
rect -34185 -88 -34045 88
rect -36405 -6320 -36265 -6130
rect -34185 -6232 -34165 -88
rect -34065 -6232 -34045 -88
rect -31875 -190 -31735 190
rect -29655 88 -29635 6232
rect -29535 88 -29515 6232
rect -27345 6130 -27205 6320
rect -25125 6232 -24985 6320
rect -29655 -88 -29515 88
rect -34185 -6320 -34045 -6232
rect -31875 -6320 -31735 -6130
rect -29655 -6232 -29635 -88
rect -29535 -6232 -29515 -88
rect -27345 -190 -27205 190
rect -25125 88 -25105 6232
rect -25005 88 -24985 6232
rect -22815 6130 -22675 6320
rect -20595 6232 -20455 6320
rect -25125 -88 -24985 88
rect -29655 -6320 -29515 -6232
rect -27345 -6320 -27205 -6130
rect -25125 -6232 -25105 -88
rect -25005 -6232 -24985 -88
rect -22815 -190 -22675 190
rect -20595 88 -20575 6232
rect -20475 88 -20455 6232
rect -18285 6130 -18145 6320
rect -16065 6232 -15925 6320
rect -20595 -88 -20455 88
rect -25125 -6320 -24985 -6232
rect -22815 -6320 -22675 -6130
rect -20595 -6232 -20575 -88
rect -20475 -6232 -20455 -88
rect -18285 -190 -18145 190
rect -16065 88 -16045 6232
rect -15945 88 -15925 6232
rect -13755 6130 -13615 6320
rect -11535 6232 -11395 6320
rect -16065 -88 -15925 88
rect -20595 -6320 -20455 -6232
rect -18285 -6320 -18145 -6130
rect -16065 -6232 -16045 -88
rect -15945 -6232 -15925 -88
rect -13755 -190 -13615 190
rect -11535 88 -11515 6232
rect -11415 88 -11395 6232
rect -9225 6130 -9085 6320
rect -7005 6232 -6865 6320
rect -11535 -88 -11395 88
rect -16065 -6320 -15925 -6232
rect -13755 -6320 -13615 -6130
rect -11535 -6232 -11515 -88
rect -11415 -6232 -11395 -88
rect -9225 -190 -9085 190
rect -7005 88 -6985 6232
rect -6885 88 -6865 6232
rect -4695 6130 -4555 6320
rect -2475 6232 -2335 6320
rect -7005 -88 -6865 88
rect -11535 -6320 -11395 -6232
rect -9225 -6320 -9085 -6130
rect -7005 -6232 -6985 -88
rect -6885 -6232 -6865 -88
rect -4695 -190 -4555 190
rect -2475 88 -2455 6232
rect -2355 88 -2335 6232
rect -165 6130 -25 6320
rect 2055 6232 2195 6320
rect -2475 -88 -2335 88
rect -7005 -6320 -6865 -6232
rect -4695 -6320 -4555 -6130
rect -2475 -6232 -2455 -88
rect -2355 -6232 -2335 -88
rect -165 -190 -25 190
rect 2055 88 2075 6232
rect 2175 88 2195 6232
rect 4365 6130 4505 6320
rect 6585 6232 6725 6320
rect 2055 -88 2195 88
rect -2475 -6320 -2335 -6232
rect -165 -6320 -25 -6130
rect 2055 -6232 2075 -88
rect 2175 -6232 2195 -88
rect 4365 -190 4505 190
rect 6585 88 6605 6232
rect 6705 88 6725 6232
rect 8895 6130 9035 6320
rect 11115 6232 11255 6320
rect 6585 -88 6725 88
rect 2055 -6320 2195 -6232
rect 4365 -6320 4505 -6130
rect 6585 -6232 6605 -88
rect 6705 -6232 6725 -88
rect 8895 -190 9035 190
rect 11115 88 11135 6232
rect 11235 88 11255 6232
rect 13425 6130 13565 6320
rect 15645 6232 15785 6320
rect 11115 -88 11255 88
rect 6585 -6320 6725 -6232
rect 8895 -6320 9035 -6130
rect 11115 -6232 11135 -88
rect 11235 -6232 11255 -88
rect 13425 -190 13565 190
rect 15645 88 15665 6232
rect 15765 88 15785 6232
rect 17955 6130 18095 6320
rect 20175 6232 20315 6320
rect 15645 -88 15785 88
rect 11115 -6320 11255 -6232
rect 13425 -6320 13565 -6130
rect 15645 -6232 15665 -88
rect 15765 -6232 15785 -88
rect 17955 -190 18095 190
rect 20175 88 20195 6232
rect 20295 88 20315 6232
rect 22485 6130 22625 6320
rect 24705 6232 24845 6320
rect 20175 -88 20315 88
rect 15645 -6320 15785 -6232
rect 17955 -6320 18095 -6130
rect 20175 -6232 20195 -88
rect 20295 -6232 20315 -88
rect 22485 -190 22625 190
rect 24705 88 24725 6232
rect 24825 88 24845 6232
rect 27015 6130 27155 6320
rect 29235 6232 29375 6320
rect 24705 -88 24845 88
rect 20175 -6320 20315 -6232
rect 22485 -6320 22625 -6130
rect 24705 -6232 24725 -88
rect 24825 -6232 24845 -88
rect 27015 -190 27155 190
rect 29235 88 29255 6232
rect 29355 88 29375 6232
rect 31545 6130 31685 6320
rect 33765 6232 33905 6320
rect 29235 -88 29375 88
rect 24705 -6320 24845 -6232
rect 27015 -6320 27155 -6130
rect 29235 -6232 29255 -88
rect 29355 -6232 29375 -88
rect 31545 -190 31685 190
rect 33765 88 33785 6232
rect 33885 88 33905 6232
rect 36075 6130 36215 6320
rect 38295 6232 38435 6320
rect 33765 -88 33905 88
rect 29235 -6320 29375 -6232
rect 31545 -6320 31685 -6130
rect 33765 -6232 33785 -88
rect 33885 -6232 33905 -88
rect 36075 -190 36215 190
rect 38295 88 38315 6232
rect 38415 88 38435 6232
rect 38295 -88 38435 88
rect 33765 -6320 33905 -6232
rect 36075 -6320 36215 -6130
rect 38295 -6232 38315 -88
rect 38415 -6232 38435 -88
rect 38295 -6320 38435 -6232
<< boundary >>
rect -38435 60 -34235 6260
rect -33905 60 -29705 6260
rect -29375 60 -25175 6260
rect -24845 60 -20645 6260
rect -20315 60 -16115 6260
rect -15785 60 -11585 6260
rect -11255 60 -7055 6260
rect -6725 60 -2525 6260
rect -2195 60 2005 6260
rect 2335 60 6535 6260
rect 6865 60 11065 6260
rect 11395 60 15595 6260
rect 15925 60 20125 6260
rect 20455 60 24655 6260
rect 24985 60 29185 6260
rect 29515 60 33715 6260
rect 34045 60 38245 6260
rect -38435 -6260 -34235 -60
rect -33905 -6260 -29705 -60
rect -29375 -6260 -25175 -60
rect -24845 -6260 -20645 -60
rect -20315 -6260 -16115 -60
rect -15785 -6260 -11585 -60
rect -11255 -6260 -7055 -60
rect -6725 -6260 -2525 -60
rect -2195 -6260 2005 -60
rect 2335 -6260 6535 -60
rect 6865 -6260 11065 -60
rect 11395 -6260 15595 -60
rect 15925 -6260 20125 -60
rect 20455 -6260 24655 -60
rect 24985 -6260 29185 -60
rect 29515 -6260 33715 -60
rect 34045 -6260 38245 -60
<< properties >>
string parameters w 20.00 l 30.00 val 617.0 carea 1.00 cperi 0.17 nx 17 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
