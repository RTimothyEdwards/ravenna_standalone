magic
tech EFXH018D
timestamp 1565723183
<< mimcap >>
rect -24830 2065 -22830 2080
rect -24830 95 -24815 2065
rect -22845 95 -22830 2065
rect -24830 80 -22830 95
rect -22565 2065 -20565 2080
rect -22565 95 -22550 2065
rect -20580 95 -20565 2065
rect -22565 80 -20565 95
rect -20300 2065 -18300 2080
rect -20300 95 -20285 2065
rect -18315 95 -18300 2065
rect -20300 80 -18300 95
rect -18035 2065 -16035 2080
rect -18035 95 -18020 2065
rect -16050 95 -16035 2065
rect -18035 80 -16035 95
rect -15770 2065 -13770 2080
rect -15770 95 -15755 2065
rect -13785 95 -13770 2065
rect -15770 80 -13770 95
rect -13505 2065 -11505 2080
rect -13505 95 -13490 2065
rect -11520 95 -11505 2065
rect -13505 80 -11505 95
rect -11240 2065 -9240 2080
rect -11240 95 -11225 2065
rect -9255 95 -9240 2065
rect -11240 80 -9240 95
rect -8975 2065 -6975 2080
rect -8975 95 -8960 2065
rect -6990 95 -6975 2065
rect -8975 80 -6975 95
rect -6710 2065 -4710 2080
rect -6710 95 -6695 2065
rect -4725 95 -4710 2065
rect -6710 80 -4710 95
rect -4445 2065 -2445 2080
rect -4445 95 -4430 2065
rect -2460 95 -2445 2065
rect -4445 80 -2445 95
rect -2180 2065 -180 2080
rect -2180 95 -2165 2065
rect -195 95 -180 2065
rect -2180 80 -180 95
rect 85 2065 2085 2080
rect 85 95 100 2065
rect 2070 95 2085 2065
rect 85 80 2085 95
rect 2350 2065 4350 2080
rect 2350 95 2365 2065
rect 4335 95 4350 2065
rect 2350 80 4350 95
rect 4615 2065 6615 2080
rect 4615 95 4630 2065
rect 6600 95 6615 2065
rect 4615 80 6615 95
rect 6880 2065 8880 2080
rect 6880 95 6895 2065
rect 8865 95 8880 2065
rect 6880 80 8880 95
rect 9145 2065 11145 2080
rect 9145 95 9160 2065
rect 11130 95 11145 2065
rect 9145 80 11145 95
rect 11410 2065 13410 2080
rect 11410 95 11425 2065
rect 13395 95 13410 2065
rect 11410 80 13410 95
rect 13675 2065 15675 2080
rect 13675 95 13690 2065
rect 15660 95 15675 2065
rect 13675 80 15675 95
rect 15940 2065 17940 2080
rect 15940 95 15955 2065
rect 17925 95 17940 2065
rect 15940 80 17940 95
rect 18205 2065 20205 2080
rect 18205 95 18220 2065
rect 20190 95 20205 2065
rect 18205 80 20205 95
rect 20470 2065 22470 2080
rect 20470 95 20485 2065
rect 22455 95 22470 2065
rect 20470 80 22470 95
rect 22735 2065 24735 2080
rect 22735 95 22750 2065
rect 24720 95 24735 2065
rect 22735 80 24735 95
rect -24830 -95 -22830 -80
rect -24830 -2065 -24815 -95
rect -22845 -2065 -22830 -95
rect -24830 -2080 -22830 -2065
rect -22565 -95 -20565 -80
rect -22565 -2065 -22550 -95
rect -20580 -2065 -20565 -95
rect -22565 -2080 -20565 -2065
rect -20300 -95 -18300 -80
rect -20300 -2065 -20285 -95
rect -18315 -2065 -18300 -95
rect -20300 -2080 -18300 -2065
rect -18035 -95 -16035 -80
rect -18035 -2065 -18020 -95
rect -16050 -2065 -16035 -95
rect -18035 -2080 -16035 -2065
rect -15770 -95 -13770 -80
rect -15770 -2065 -15755 -95
rect -13785 -2065 -13770 -95
rect -15770 -2080 -13770 -2065
rect -13505 -95 -11505 -80
rect -13505 -2065 -13490 -95
rect -11520 -2065 -11505 -95
rect -13505 -2080 -11505 -2065
rect -11240 -95 -9240 -80
rect -11240 -2065 -11225 -95
rect -9255 -2065 -9240 -95
rect -11240 -2080 -9240 -2065
rect -8975 -95 -6975 -80
rect -8975 -2065 -8960 -95
rect -6990 -2065 -6975 -95
rect -8975 -2080 -6975 -2065
rect -6710 -95 -4710 -80
rect -6710 -2065 -6695 -95
rect -4725 -2065 -4710 -95
rect -6710 -2080 -4710 -2065
rect -4445 -95 -2445 -80
rect -4445 -2065 -4430 -95
rect -2460 -2065 -2445 -95
rect -4445 -2080 -2445 -2065
rect -2180 -95 -180 -80
rect -2180 -2065 -2165 -95
rect -195 -2065 -180 -95
rect -2180 -2080 -180 -2065
rect 85 -95 2085 -80
rect 85 -2065 100 -95
rect 2070 -2065 2085 -95
rect 85 -2080 2085 -2065
rect 2350 -95 4350 -80
rect 2350 -2065 2365 -95
rect 4335 -2065 4350 -95
rect 2350 -2080 4350 -2065
rect 4615 -95 6615 -80
rect 4615 -2065 4630 -95
rect 6600 -2065 6615 -95
rect 4615 -2080 6615 -2065
rect 6880 -95 8880 -80
rect 6880 -2065 6895 -95
rect 8865 -2065 8880 -95
rect 6880 -2080 8880 -2065
rect 9145 -95 11145 -80
rect 9145 -2065 9160 -95
rect 11130 -2065 11145 -95
rect 9145 -2080 11145 -2065
rect 11410 -95 13410 -80
rect 11410 -2065 11425 -95
rect 13395 -2065 13410 -95
rect 11410 -2080 13410 -2065
rect 13675 -95 15675 -80
rect 13675 -2065 13690 -95
rect 15660 -2065 15675 -95
rect 13675 -2080 15675 -2065
rect 15940 -95 17940 -80
rect 15940 -2065 15955 -95
rect 17925 -2065 17940 -95
rect 15940 -2080 17940 -2065
rect 18205 -95 20205 -80
rect 18205 -2065 18220 -95
rect 20190 -2065 20205 -95
rect 18205 -2080 20205 -2065
rect 20470 -95 22470 -80
rect 20470 -2065 20485 -95
rect 22455 -2065 22470 -95
rect 20470 -2080 22470 -2065
rect 22735 -95 24735 -80
rect 22735 -2065 22750 -95
rect 24720 -2065 24735 -95
rect 22735 -2080 24735 -2065
<< mimcapcontact >>
rect -24815 95 -22845 2065
rect -22550 95 -20580 2065
rect -20285 95 -18315 2065
rect -18020 95 -16050 2065
rect -15755 95 -13785 2065
rect -13490 95 -11520 2065
rect -11225 95 -9255 2065
rect -8960 95 -6990 2065
rect -6695 95 -4725 2065
rect -4430 95 -2460 2065
rect -2165 95 -195 2065
rect 100 95 2070 2065
rect 2365 95 4335 2065
rect 4630 95 6600 2065
rect 6895 95 8865 2065
rect 9160 95 11130 2065
rect 11425 95 13395 2065
rect 13690 95 15660 2065
rect 15955 95 17925 2065
rect 18220 95 20190 2065
rect 20485 95 22455 2065
rect 22750 95 24720 2065
rect -24815 -2065 -22845 -95
rect -22550 -2065 -20580 -95
rect -20285 -2065 -18315 -95
rect -18020 -2065 -16050 -95
rect -15755 -2065 -13785 -95
rect -13490 -2065 -11520 -95
rect -11225 -2065 -9255 -95
rect -8960 -2065 -6990 -95
rect -6695 -2065 -4725 -95
rect -4430 -2065 -2460 -95
rect -2165 -2065 -195 -95
rect 100 -2065 2070 -95
rect 2365 -2065 4335 -95
rect 4630 -2065 6600 -95
rect 6895 -2065 8865 -95
rect 9160 -2065 11130 -95
rect 11425 -2065 13395 -95
rect 13690 -2065 15660 -95
rect 15955 -2065 17925 -95
rect 18220 -2065 20190 -95
rect 20485 -2065 22455 -95
rect 22750 -2065 24720 -95
<< metal4 >>
rect -24880 2116 -22685 2130
rect -24880 2080 -22745 2116
rect -24880 80 -24830 2080
rect -22830 80 -22745 2080
rect -24880 44 -22745 80
rect -22695 44 -22685 2116
rect -24880 30 -22685 44
rect -22615 2116 -20420 2130
rect -22615 2080 -20480 2116
rect -22615 80 -22565 2080
rect -20565 80 -20480 2080
rect -22615 44 -20480 80
rect -20430 44 -20420 2116
rect -22615 30 -20420 44
rect -20350 2116 -18155 2130
rect -20350 2080 -18215 2116
rect -20350 80 -20300 2080
rect -18300 80 -18215 2080
rect -20350 44 -18215 80
rect -18165 44 -18155 2116
rect -20350 30 -18155 44
rect -18085 2116 -15890 2130
rect -18085 2080 -15950 2116
rect -18085 80 -18035 2080
rect -16035 80 -15950 2080
rect -18085 44 -15950 80
rect -15900 44 -15890 2116
rect -18085 30 -15890 44
rect -15820 2116 -13625 2130
rect -15820 2080 -13685 2116
rect -15820 80 -15770 2080
rect -13770 80 -13685 2080
rect -15820 44 -13685 80
rect -13635 44 -13625 2116
rect -15820 30 -13625 44
rect -13555 2116 -11360 2130
rect -13555 2080 -11420 2116
rect -13555 80 -13505 2080
rect -11505 80 -11420 2080
rect -13555 44 -11420 80
rect -11370 44 -11360 2116
rect -13555 30 -11360 44
rect -11290 2116 -9095 2130
rect -11290 2080 -9155 2116
rect -11290 80 -11240 2080
rect -9240 80 -9155 2080
rect -11290 44 -9155 80
rect -9105 44 -9095 2116
rect -11290 30 -9095 44
rect -9025 2116 -6830 2130
rect -9025 2080 -6890 2116
rect -9025 80 -8975 2080
rect -6975 80 -6890 2080
rect -9025 44 -6890 80
rect -6840 44 -6830 2116
rect -9025 30 -6830 44
rect -6760 2116 -4565 2130
rect -6760 2080 -4625 2116
rect -6760 80 -6710 2080
rect -4710 80 -4625 2080
rect -6760 44 -4625 80
rect -4575 44 -4565 2116
rect -6760 30 -4565 44
rect -4495 2116 -2300 2130
rect -4495 2080 -2360 2116
rect -4495 80 -4445 2080
rect -2445 80 -2360 2080
rect -4495 44 -2360 80
rect -2310 44 -2300 2116
rect -4495 30 -2300 44
rect -2230 2116 -35 2130
rect -2230 2080 -95 2116
rect -2230 80 -2180 2080
rect -180 80 -95 2080
rect -2230 44 -95 80
rect -45 44 -35 2116
rect -2230 30 -35 44
rect 35 2116 2230 2130
rect 35 2080 2170 2116
rect 35 80 85 2080
rect 2085 80 2170 2080
rect 35 44 2170 80
rect 2220 44 2230 2116
rect 35 30 2230 44
rect 2300 2116 4495 2130
rect 2300 2080 4435 2116
rect 2300 80 2350 2080
rect 4350 80 4435 2080
rect 2300 44 4435 80
rect 4485 44 4495 2116
rect 2300 30 4495 44
rect 4565 2116 6760 2130
rect 4565 2080 6700 2116
rect 4565 80 4615 2080
rect 6615 80 6700 2080
rect 4565 44 6700 80
rect 6750 44 6760 2116
rect 4565 30 6760 44
rect 6830 2116 9025 2130
rect 6830 2080 8965 2116
rect 6830 80 6880 2080
rect 8880 80 8965 2080
rect 6830 44 8965 80
rect 9015 44 9025 2116
rect 6830 30 9025 44
rect 9095 2116 11290 2130
rect 9095 2080 11230 2116
rect 9095 80 9145 2080
rect 11145 80 11230 2080
rect 9095 44 11230 80
rect 11280 44 11290 2116
rect 9095 30 11290 44
rect 11360 2116 13555 2130
rect 11360 2080 13495 2116
rect 11360 80 11410 2080
rect 13410 80 13495 2080
rect 11360 44 13495 80
rect 13545 44 13555 2116
rect 11360 30 13555 44
rect 13625 2116 15820 2130
rect 13625 2080 15760 2116
rect 13625 80 13675 2080
rect 15675 80 15760 2080
rect 13625 44 15760 80
rect 15810 44 15820 2116
rect 13625 30 15820 44
rect 15890 2116 18085 2130
rect 15890 2080 18025 2116
rect 15890 80 15940 2080
rect 17940 80 18025 2080
rect 15890 44 18025 80
rect 18075 44 18085 2116
rect 15890 30 18085 44
rect 18155 2116 20350 2130
rect 18155 2080 20290 2116
rect 18155 80 18205 2080
rect 20205 80 20290 2080
rect 18155 44 20290 80
rect 20340 44 20350 2116
rect 18155 30 20350 44
rect 20420 2116 22615 2130
rect 20420 2080 22555 2116
rect 20420 80 20470 2080
rect 22470 80 22555 2080
rect 20420 44 22555 80
rect 22605 44 22615 2116
rect 20420 30 22615 44
rect 22685 2116 24880 2130
rect 22685 2080 24820 2116
rect 22685 80 22735 2080
rect 24735 80 24820 2080
rect 22685 44 24820 80
rect 24870 44 24880 2116
rect 22685 30 24880 44
rect -24880 -44 -22685 -30
rect -24880 -80 -22745 -44
rect -24880 -2080 -24830 -80
rect -22830 -2080 -22745 -80
rect -24880 -2116 -22745 -2080
rect -22695 -2116 -22685 -44
rect -24880 -2130 -22685 -2116
rect -22615 -44 -20420 -30
rect -22615 -80 -20480 -44
rect -22615 -2080 -22565 -80
rect -20565 -2080 -20480 -80
rect -22615 -2116 -20480 -2080
rect -20430 -2116 -20420 -44
rect -22615 -2130 -20420 -2116
rect -20350 -44 -18155 -30
rect -20350 -80 -18215 -44
rect -20350 -2080 -20300 -80
rect -18300 -2080 -18215 -80
rect -20350 -2116 -18215 -2080
rect -18165 -2116 -18155 -44
rect -20350 -2130 -18155 -2116
rect -18085 -44 -15890 -30
rect -18085 -80 -15950 -44
rect -18085 -2080 -18035 -80
rect -16035 -2080 -15950 -80
rect -18085 -2116 -15950 -2080
rect -15900 -2116 -15890 -44
rect -18085 -2130 -15890 -2116
rect -15820 -44 -13625 -30
rect -15820 -80 -13685 -44
rect -15820 -2080 -15770 -80
rect -13770 -2080 -13685 -80
rect -15820 -2116 -13685 -2080
rect -13635 -2116 -13625 -44
rect -15820 -2130 -13625 -2116
rect -13555 -44 -11360 -30
rect -13555 -80 -11420 -44
rect -13555 -2080 -13505 -80
rect -11505 -2080 -11420 -80
rect -13555 -2116 -11420 -2080
rect -11370 -2116 -11360 -44
rect -13555 -2130 -11360 -2116
rect -11290 -44 -9095 -30
rect -11290 -80 -9155 -44
rect -11290 -2080 -11240 -80
rect -9240 -2080 -9155 -80
rect -11290 -2116 -9155 -2080
rect -9105 -2116 -9095 -44
rect -11290 -2130 -9095 -2116
rect -9025 -44 -6830 -30
rect -9025 -80 -6890 -44
rect -9025 -2080 -8975 -80
rect -6975 -2080 -6890 -80
rect -9025 -2116 -6890 -2080
rect -6840 -2116 -6830 -44
rect -9025 -2130 -6830 -2116
rect -6760 -44 -4565 -30
rect -6760 -80 -4625 -44
rect -6760 -2080 -6710 -80
rect -4710 -2080 -4625 -80
rect -6760 -2116 -4625 -2080
rect -4575 -2116 -4565 -44
rect -6760 -2130 -4565 -2116
rect -4495 -44 -2300 -30
rect -4495 -80 -2360 -44
rect -4495 -2080 -4445 -80
rect -2445 -2080 -2360 -80
rect -4495 -2116 -2360 -2080
rect -2310 -2116 -2300 -44
rect -4495 -2130 -2300 -2116
rect -2230 -44 -35 -30
rect -2230 -80 -95 -44
rect -2230 -2080 -2180 -80
rect -180 -2080 -95 -80
rect -2230 -2116 -95 -2080
rect -45 -2116 -35 -44
rect -2230 -2130 -35 -2116
rect 35 -44 2230 -30
rect 35 -80 2170 -44
rect 35 -2080 85 -80
rect 2085 -2080 2170 -80
rect 35 -2116 2170 -2080
rect 2220 -2116 2230 -44
rect 35 -2130 2230 -2116
rect 2300 -44 4495 -30
rect 2300 -80 4435 -44
rect 2300 -2080 2350 -80
rect 4350 -2080 4435 -80
rect 2300 -2116 4435 -2080
rect 4485 -2116 4495 -44
rect 2300 -2130 4495 -2116
rect 4565 -44 6760 -30
rect 4565 -80 6700 -44
rect 4565 -2080 4615 -80
rect 6615 -2080 6700 -80
rect 4565 -2116 6700 -2080
rect 6750 -2116 6760 -44
rect 4565 -2130 6760 -2116
rect 6830 -44 9025 -30
rect 6830 -80 8965 -44
rect 6830 -2080 6880 -80
rect 8880 -2080 8965 -80
rect 6830 -2116 8965 -2080
rect 9015 -2116 9025 -44
rect 6830 -2130 9025 -2116
rect 9095 -44 11290 -30
rect 9095 -80 11230 -44
rect 9095 -2080 9145 -80
rect 11145 -2080 11230 -80
rect 9095 -2116 11230 -2080
rect 11280 -2116 11290 -44
rect 9095 -2130 11290 -2116
rect 11360 -44 13555 -30
rect 11360 -80 13495 -44
rect 11360 -2080 11410 -80
rect 13410 -2080 13495 -80
rect 11360 -2116 13495 -2080
rect 13545 -2116 13555 -44
rect 11360 -2130 13555 -2116
rect 13625 -44 15820 -30
rect 13625 -80 15760 -44
rect 13625 -2080 13675 -80
rect 15675 -2080 15760 -80
rect 13625 -2116 15760 -2080
rect 15810 -2116 15820 -44
rect 13625 -2130 15820 -2116
rect 15890 -44 18085 -30
rect 15890 -80 18025 -44
rect 15890 -2080 15940 -80
rect 17940 -2080 18025 -80
rect 15890 -2116 18025 -2080
rect 18075 -2116 18085 -44
rect 15890 -2130 18085 -2116
rect 18155 -44 20350 -30
rect 18155 -80 20290 -44
rect 18155 -2080 18205 -80
rect 20205 -2080 20290 -80
rect 18155 -2116 20290 -2080
rect 20340 -2116 20350 -44
rect 18155 -2130 20350 -2116
rect 20420 -44 22615 -30
rect 20420 -80 22555 -44
rect 20420 -2080 20470 -80
rect 22470 -2080 22555 -80
rect 20420 -2116 22555 -2080
rect 22605 -2116 22615 -44
rect 20420 -2130 22615 -2116
rect 22685 -44 24880 -30
rect 22685 -80 24820 -44
rect 22685 -2080 22735 -80
rect 24735 -2080 24820 -80
rect 22685 -2116 24820 -2080
rect 24870 -2116 24880 -44
rect 22685 -2130 24880 -2116
<< viatp >>
rect -22745 44 -22695 2116
rect -20480 44 -20430 2116
rect -18215 44 -18165 2116
rect -15950 44 -15900 2116
rect -13685 44 -13635 2116
rect -11420 44 -11370 2116
rect -9155 44 -9105 2116
rect -6890 44 -6840 2116
rect -4625 44 -4575 2116
rect -2360 44 -2310 2116
rect -95 44 -45 2116
rect 2170 44 2220 2116
rect 4435 44 4485 2116
rect 6700 44 6750 2116
rect 8965 44 9015 2116
rect 11230 44 11280 2116
rect 13495 44 13545 2116
rect 15760 44 15810 2116
rect 18025 44 18075 2116
rect 20290 44 20340 2116
rect 22555 44 22605 2116
rect 24820 44 24870 2116
rect -22745 -2116 -22695 -44
rect -20480 -2116 -20430 -44
rect -18215 -2116 -18165 -44
rect -15950 -2116 -15900 -44
rect -13685 -2116 -13635 -44
rect -11420 -2116 -11370 -44
rect -9155 -2116 -9105 -44
rect -6890 -2116 -6840 -44
rect -4625 -2116 -4575 -44
rect -2360 -2116 -2310 -44
rect -95 -2116 -45 -44
rect 2170 -2116 2220 -44
rect 4435 -2116 4485 -44
rect 6700 -2116 6750 -44
rect 8965 -2116 9015 -44
rect 11230 -2116 11280 -44
rect 13495 -2116 13545 -44
rect 15760 -2116 15810 -44
rect 18025 -2116 18075 -44
rect 20290 -2116 20340 -44
rect 22555 -2116 22605 -44
rect 24820 -2116 24870 -44
<< metaltp >>
rect -23865 2065 -23795 2160
rect -22755 2116 -22685 2160
rect -23865 -95 -23795 95
rect -22755 44 -22745 2116
rect -22695 44 -22685 2116
rect -21600 2065 -21530 2160
rect -20490 2116 -20420 2160
rect -22755 -44 -22685 44
rect -23865 -2160 -23795 -2065
rect -22755 -2116 -22745 -44
rect -22695 -2116 -22685 -44
rect -21600 -95 -21530 95
rect -20490 44 -20480 2116
rect -20430 44 -20420 2116
rect -19335 2065 -19265 2160
rect -18225 2116 -18155 2160
rect -20490 -44 -20420 44
rect -22755 -2160 -22685 -2116
rect -21600 -2160 -21530 -2065
rect -20490 -2116 -20480 -44
rect -20430 -2116 -20420 -44
rect -19335 -95 -19265 95
rect -18225 44 -18215 2116
rect -18165 44 -18155 2116
rect -17070 2065 -17000 2160
rect -15960 2116 -15890 2160
rect -18225 -44 -18155 44
rect -20490 -2160 -20420 -2116
rect -19335 -2160 -19265 -2065
rect -18225 -2116 -18215 -44
rect -18165 -2116 -18155 -44
rect -17070 -95 -17000 95
rect -15960 44 -15950 2116
rect -15900 44 -15890 2116
rect -14805 2065 -14735 2160
rect -13695 2116 -13625 2160
rect -15960 -44 -15890 44
rect -18225 -2160 -18155 -2116
rect -17070 -2160 -17000 -2065
rect -15960 -2116 -15950 -44
rect -15900 -2116 -15890 -44
rect -14805 -95 -14735 95
rect -13695 44 -13685 2116
rect -13635 44 -13625 2116
rect -12540 2065 -12470 2160
rect -11430 2116 -11360 2160
rect -13695 -44 -13625 44
rect -15960 -2160 -15890 -2116
rect -14805 -2160 -14735 -2065
rect -13695 -2116 -13685 -44
rect -13635 -2116 -13625 -44
rect -12540 -95 -12470 95
rect -11430 44 -11420 2116
rect -11370 44 -11360 2116
rect -10275 2065 -10205 2160
rect -9165 2116 -9095 2160
rect -11430 -44 -11360 44
rect -13695 -2160 -13625 -2116
rect -12540 -2160 -12470 -2065
rect -11430 -2116 -11420 -44
rect -11370 -2116 -11360 -44
rect -10275 -95 -10205 95
rect -9165 44 -9155 2116
rect -9105 44 -9095 2116
rect -8010 2065 -7940 2160
rect -6900 2116 -6830 2160
rect -9165 -44 -9095 44
rect -11430 -2160 -11360 -2116
rect -10275 -2160 -10205 -2065
rect -9165 -2116 -9155 -44
rect -9105 -2116 -9095 -44
rect -8010 -95 -7940 95
rect -6900 44 -6890 2116
rect -6840 44 -6830 2116
rect -5745 2065 -5675 2160
rect -4635 2116 -4565 2160
rect -6900 -44 -6830 44
rect -9165 -2160 -9095 -2116
rect -8010 -2160 -7940 -2065
rect -6900 -2116 -6890 -44
rect -6840 -2116 -6830 -44
rect -5745 -95 -5675 95
rect -4635 44 -4625 2116
rect -4575 44 -4565 2116
rect -3480 2065 -3410 2160
rect -2370 2116 -2300 2160
rect -4635 -44 -4565 44
rect -6900 -2160 -6830 -2116
rect -5745 -2160 -5675 -2065
rect -4635 -2116 -4625 -44
rect -4575 -2116 -4565 -44
rect -3480 -95 -3410 95
rect -2370 44 -2360 2116
rect -2310 44 -2300 2116
rect -1215 2065 -1145 2160
rect -105 2116 -35 2160
rect -2370 -44 -2300 44
rect -4635 -2160 -4565 -2116
rect -3480 -2160 -3410 -2065
rect -2370 -2116 -2360 -44
rect -2310 -2116 -2300 -44
rect -1215 -95 -1145 95
rect -105 44 -95 2116
rect -45 44 -35 2116
rect 1050 2065 1120 2160
rect 2160 2116 2230 2160
rect -105 -44 -35 44
rect -2370 -2160 -2300 -2116
rect -1215 -2160 -1145 -2065
rect -105 -2116 -95 -44
rect -45 -2116 -35 -44
rect 1050 -95 1120 95
rect 2160 44 2170 2116
rect 2220 44 2230 2116
rect 3315 2065 3385 2160
rect 4425 2116 4495 2160
rect 2160 -44 2230 44
rect -105 -2160 -35 -2116
rect 1050 -2160 1120 -2065
rect 2160 -2116 2170 -44
rect 2220 -2116 2230 -44
rect 3315 -95 3385 95
rect 4425 44 4435 2116
rect 4485 44 4495 2116
rect 5580 2065 5650 2160
rect 6690 2116 6760 2160
rect 4425 -44 4495 44
rect 2160 -2160 2230 -2116
rect 3315 -2160 3385 -2065
rect 4425 -2116 4435 -44
rect 4485 -2116 4495 -44
rect 5580 -95 5650 95
rect 6690 44 6700 2116
rect 6750 44 6760 2116
rect 7845 2065 7915 2160
rect 8955 2116 9025 2160
rect 6690 -44 6760 44
rect 4425 -2160 4495 -2116
rect 5580 -2160 5650 -2065
rect 6690 -2116 6700 -44
rect 6750 -2116 6760 -44
rect 7845 -95 7915 95
rect 8955 44 8965 2116
rect 9015 44 9025 2116
rect 10110 2065 10180 2160
rect 11220 2116 11290 2160
rect 8955 -44 9025 44
rect 6690 -2160 6760 -2116
rect 7845 -2160 7915 -2065
rect 8955 -2116 8965 -44
rect 9015 -2116 9025 -44
rect 10110 -95 10180 95
rect 11220 44 11230 2116
rect 11280 44 11290 2116
rect 12375 2065 12445 2160
rect 13485 2116 13555 2160
rect 11220 -44 11290 44
rect 8955 -2160 9025 -2116
rect 10110 -2160 10180 -2065
rect 11220 -2116 11230 -44
rect 11280 -2116 11290 -44
rect 12375 -95 12445 95
rect 13485 44 13495 2116
rect 13545 44 13555 2116
rect 14640 2065 14710 2160
rect 15750 2116 15820 2160
rect 13485 -44 13555 44
rect 11220 -2160 11290 -2116
rect 12375 -2160 12445 -2065
rect 13485 -2116 13495 -44
rect 13545 -2116 13555 -44
rect 14640 -95 14710 95
rect 15750 44 15760 2116
rect 15810 44 15820 2116
rect 16905 2065 16975 2160
rect 18015 2116 18085 2160
rect 15750 -44 15820 44
rect 13485 -2160 13555 -2116
rect 14640 -2160 14710 -2065
rect 15750 -2116 15760 -44
rect 15810 -2116 15820 -44
rect 16905 -95 16975 95
rect 18015 44 18025 2116
rect 18075 44 18085 2116
rect 19170 2065 19240 2160
rect 20280 2116 20350 2160
rect 18015 -44 18085 44
rect 15750 -2160 15820 -2116
rect 16905 -2160 16975 -2065
rect 18015 -2116 18025 -44
rect 18075 -2116 18085 -44
rect 19170 -95 19240 95
rect 20280 44 20290 2116
rect 20340 44 20350 2116
rect 21435 2065 21505 2160
rect 22545 2116 22615 2160
rect 20280 -44 20350 44
rect 18015 -2160 18085 -2116
rect 19170 -2160 19240 -2065
rect 20280 -2116 20290 -44
rect 20340 -2116 20350 -44
rect 21435 -95 21505 95
rect 22545 44 22555 2116
rect 22605 44 22615 2116
rect 23700 2065 23770 2160
rect 24810 2116 24880 2160
rect 22545 -44 22615 44
rect 20280 -2160 20350 -2116
rect 21435 -2160 21505 -2065
rect 22545 -2116 22555 -44
rect 22605 -2116 22615 -44
rect 23700 -95 23770 95
rect 24810 44 24820 2116
rect 24870 44 24880 2116
rect 24810 -44 24880 44
rect 22545 -2160 22615 -2116
rect 23700 -2160 23770 -2065
rect 24810 -2116 24820 -44
rect 24870 -2116 24880 -44
rect 24810 -2160 24880 -2116
<< properties >>
string parameters w 20.00 l 20.00 val 413.6 carea 1.00 cperi 0.17 nx 22 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
