magic
tech EFXH018D
timestamp 1494891594
<< metal2 >>
rect 0 96 96 960
rect 0 0 528 96
<< end >>
