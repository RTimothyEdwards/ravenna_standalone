magic
tech EFXH018A
magscale 1 2
timestamp 1527118791
<< checkpaint >>
rect 3982 -3710 13512 4880
<< metal1 >>
rect 6034 2580 6234 2880
rect 6064 2578 6134 2580
rect 7174 2530 7374 2870
rect 7908 2576 8108 2878
rect 8648 2576 8848 2876
rect 9384 2576 9584 2878
rect 11258 2578 11458 2880
rect 6094 2424 11468 2530
rect 6094 2268 6140 2424
rect 6780 2268 6826 2424
rect 7260 2268 7306 2424
rect 7760 2268 7806 2424
rect 6094 1846 6144 2268
rect 6240 2224 6288 2246
rect 6096 1840 6144 1846
rect 6238 1862 6288 2224
rect 6636 2230 6684 2246
rect 6636 1862 6686 2230
rect 6238 1596 6284 1862
rect 6050 1508 6284 1596
rect 6100 1278 6148 1280
rect 6092 852 6148 1278
rect 6238 1258 6284 1508
rect 6640 1258 6686 1862
rect 6780 1840 6828 2268
rect 7122 2238 7170 2246
rect 7122 1862 7180 2238
rect 6784 1270 6832 1280
rect 6238 874 6292 1258
rect 6640 1094 6688 1258
rect 6776 1094 6832 1270
rect 6640 978 6832 1094
rect 6640 874 6688 978
rect 6238 872 6284 874
rect 6640 864 6686 874
rect 6776 852 6832 978
rect 7134 1738 7180 1862
rect 7260 1842 7314 2268
rect 7410 1862 7458 2246
rect 7266 1840 7314 1842
rect 7412 1738 7458 1862
rect 7134 1480 7476 1738
rect 7752 1844 7806 2268
rect 7896 1862 7944 2246
rect 8292 2234 8340 2246
rect 8292 2124 8344 2234
rect 8292 1972 8358 2124
rect 8292 1862 8344 1972
rect 7752 1840 7800 1844
rect 7134 1258 7180 1480
rect 7126 876 7180 1258
rect 7126 874 7174 876
rect 7270 852 7318 1280
rect 7412 1258 7458 1480
rect 7756 1266 7804 1280
rect 7412 874 7462 1258
rect 7752 1122 7804 1266
rect 7896 1258 7942 1862
rect 8298 1258 8344 1862
rect 8436 1794 8514 2424
rect 7896 1122 7948 1258
rect 7752 1024 7948 1122
rect 7412 868 7458 874
rect 7752 852 7804 1024
rect 7896 874 7948 1024
rect 8296 874 8344 1258
rect 7896 870 7942 874
rect 8298 868 8344 874
rect 8440 1264 8488 1280
rect 8440 852 8490 1264
rect 6092 696 6146 852
rect 6776 696 6822 852
rect 7270 696 7316 852
rect 7752 696 7798 852
rect 8444 696 8490 852
rect 8680 786 8822 2424
rect 8976 2268 9052 2424
rect 9690 2268 9736 2424
rect 10186 2268 10232 2424
rect 10672 2268 10718 2424
rect 8976 1840 9066 2268
rect 9162 2124 9210 2246
rect 9146 1972 9210 2124
rect 9162 1862 9210 1972
rect 9558 2234 9606 2246
rect 9556 1862 9606 2234
rect 8976 1794 9052 1840
rect 9014 852 9062 1280
rect 9162 1258 9208 1862
rect 9158 874 9208 1258
rect 9556 1258 9602 1862
rect 9690 1844 9750 2268
rect 9702 1840 9750 1844
rect 10044 1862 10092 2246
rect 10044 1738 10090 1862
rect 10186 1842 10236 2268
rect 10332 2238 10380 2246
rect 10188 1840 10236 1842
rect 10330 1862 10380 2238
rect 10330 1738 10376 1862
rect 9554 1122 9602 1258
rect 9698 1122 9746 1280
rect 9958 1480 10376 1738
rect 10044 1258 10090 1480
rect 9554 1024 9746 1122
rect 9554 874 9602 1024
rect 9162 868 9208 874
rect 9556 870 9602 874
rect 9016 696 9062 852
rect 9698 852 9746 1024
rect 10040 874 10090 1258
rect 10044 868 10090 874
rect 10184 1260 10232 1280
rect 10184 852 10240 1260
rect 10330 1258 10376 1480
rect 10672 1842 10722 2268
rect 10818 1862 10866 2246
rect 10674 1840 10722 1842
rect 10328 874 10376 1258
rect 10670 1270 10718 1280
rect 10670 1094 10722 1270
rect 10820 1258 10866 1862
rect 11214 2224 11262 2246
rect 11212 1862 11262 2224
rect 10814 1094 10866 1258
rect 10670 978 10866 1094
rect 10670 852 10722 978
rect 10814 874 10866 978
rect 11212 1666 11258 1862
rect 11358 1852 11468 2424
rect 11358 1840 11406 1852
rect 11212 1498 11442 1666
rect 11212 1258 11258 1498
rect 11210 874 11258 1258
rect 11354 1266 11402 1280
rect 10820 864 10866 874
rect 11354 852 11464 1266
rect 9698 696 9744 852
rect 10194 696 10240 852
rect 10676 696 10722 852
rect 11358 696 11464 852
rect 5994 592 11464 696
rect 5994 546 6516 592
rect 7998 546 8164 592
rect 9330 546 9494 592
rect 10962 590 11464 592
rect 10962 546 11216 590
rect 5994 386 11216 546
rect 5994 384 6324 386
rect 5986 -34 6186 46
rect 5986 -154 6280 -34
rect 8678 -234 8826 226
rect 8716 -350 8788 -234
rect 6288 -510 11216 -350
rect 6528 -606 6744 -510
rect 8678 -606 8826 -510
rect 10760 -606 10976 -510
rect 6272 -766 11232 -606
rect 5988 -986 6188 -886
rect 5988 -1086 6292 -986
rect 6762 -974 6828 -766
rect 7128 -866 7208 -766
rect 7516 -884 7582 -766
rect 7860 -884 7956 -838
rect 5982 -1394 6365 -1194
rect 7910 -932 7956 -884
rect 8016 -886 9488 -812
rect 9548 -884 9644 -838
rect 9922 -884 9988 -766
rect 10296 -866 10376 -766
rect 7910 -978 8220 -932
rect 8266 -936 9238 -886
rect 9548 -932 9594 -884
rect 6760 -1502 6824 -1326
rect 7134 -1502 7204 -1374
rect 7514 -1502 7584 -1344
rect 8156 -1058 8220 -978
rect 8156 -1114 8350 -1058
rect 8246 -1142 8350 -1114
rect 8246 -1228 8380 -1142
rect 7882 -1502 7968 -1382
rect 8222 -1502 8286 -1366
rect 8676 -1420 8832 -936
rect 9284 -978 9594 -932
rect 9284 -1058 9348 -978
rect 9154 -1114 9348 -1058
rect 9154 -1142 9258 -1114
rect 9124 -1228 9258 -1142
rect 10676 -974 10742 -766
rect 9218 -1502 9282 -1366
rect 9536 -1502 9622 -1382
rect 9920 -1502 9990 -1344
rect 10300 -1502 10370 -1374
rect 10680 -1502 10744 -1326
rect 11304 -1502 11464 590
rect 6272 -1662 11464 -1502
rect 11304 -1664 11464 -1662
<< obsm1 >>
rect 6328 2358 6400 2378
rect 6526 2360 6598 2378
rect 6302 2292 6432 2358
rect 6500 2292 6630 2360
rect 7012 2358 7084 2378
rect 6990 2292 7120 2358
rect 7498 2360 7570 2378
rect 7468 2292 7596 2360
rect 7984 2358 8056 2378
rect 8182 2360 8254 2378
rect 7950 2292 8080 2358
rect 8148 2292 8276 2360
rect 6438 2228 6486 2246
rect 6438 1862 6488 2228
rect 6440 1666 6488 1862
rect 6336 1510 6590 1666
rect 6440 1258 6488 1510
rect 6924 2232 6972 2246
rect 6924 1862 6974 2232
rect 6928 1604 6974 1862
rect 6844 1504 6974 1604
rect 6440 888 6490 1258
rect 6442 874 6490 888
rect 6928 1258 6974 1504
rect 7608 1862 7656 2246
rect 7610 1604 7656 1862
rect 8094 2232 8142 2246
rect 8092 1862 8142 2232
rect 7610 1504 7758 1604
rect 6928 874 6976 1258
rect 7610 1258 7656 1504
rect 7610 874 7660 1258
rect 8092 1668 8140 1862
rect 7988 1510 8244 1668
rect 8092 1258 8140 1510
rect 7610 872 7656 874
rect 8092 892 8146 1258
rect 8098 874 8146 892
rect 6302 744 6436 810
rect 6502 744 6634 810
rect 6332 742 6404 744
rect 6530 742 6602 744
rect 6986 744 7120 810
rect 7016 742 7088 744
rect 7474 744 7606 810
rect 7502 742 7574 744
rect 7958 744 8092 810
rect 8162 744 8294 810
rect 7988 742 8060 744
rect 8186 742 8258 744
rect 9250 2360 9322 2378
rect 9222 2292 9350 2360
rect 9448 2358 9520 2378
rect 9418 2292 9548 2358
rect 9934 2360 10006 2378
rect 9906 2292 10034 2360
rect 10420 2358 10492 2378
rect 10390 2292 10520 2358
rect 10906 2360 10978 2378
rect 10874 2292 11006 2360
rect 11104 2358 11176 2378
rect 11074 2292 11204 2358
rect 9360 2244 9408 2246
rect 9354 1862 9408 2244
rect 9260 1668 9306 1678
rect 9354 1668 9404 1862
rect 9460 1668 9506 1678
rect 9260 1510 9506 1668
rect 9260 1500 9306 1510
rect 9354 884 9404 1510
rect 9460 1500 9506 1510
rect 9846 1862 9894 2246
rect 9848 1604 9894 1862
rect 10530 2232 10578 2246
rect 10528 1862 10578 2232
rect 9746 1504 9894 1604
rect 9356 874 9404 884
rect 9848 1258 9894 1504
rect 9842 874 9894 1258
rect 9848 872 9894 874
rect 10528 1604 10574 1862
rect 11016 2242 11064 2246
rect 10528 1504 10684 1604
rect 10528 1258 10574 1504
rect 10526 874 10574 1258
rect 10912 1666 10958 1678
rect 11012 1666 11064 2242
rect 11114 1666 11160 1678
rect 10912 1508 11160 1666
rect 10912 1500 10958 1508
rect 11012 878 11064 1508
rect 11114 1500 11160 1508
rect 11012 874 11060 878
rect 9220 744 9350 810
rect 9418 744 9552 810
rect 9246 742 9318 744
rect 9444 742 9516 744
rect 9900 744 10030 810
rect 9930 742 10002 744
rect 10386 744 10520 810
rect 10416 742 10488 744
rect 10872 744 11002 810
rect 11070 744 11204 810
rect 10902 742 10974 744
rect 11100 742 11172 744
rect 6324 324 6382 386
rect 6642 324 6700 386
rect 6772 270 6830 386
rect 6876 270 7380 326
rect 7426 270 7484 386
rect 7556 270 7614 386
rect 7660 270 8164 326
rect 8210 270 8268 386
rect 8340 324 8398 386
rect 8658 324 8716 386
rect 8788 324 8846 386
rect 9106 324 9164 386
rect 9236 270 9294 386
rect 9340 270 9844 326
rect 9890 270 9948 386
rect 10020 270 10078 386
rect 10124 270 10628 326
rect 10674 270 10732 386
rect 10804 324 10862 386
rect 11122 324 11180 386
rect 6428 164 6790 222
rect 6428 -23 6484 164
rect 6540 36 6770 112
rect 6876 40 6942 270
rect 6988 112 7044 220
rect 7094 158 7268 224
rect 6988 36 7166 112
rect 6708 -10 6770 36
rect 7212 -10 7268 158
rect 7314 96 7380 270
rect 7660 96 7726 270
rect 7314 40 7486 96
rect 6428 -85 6544 -23
rect 6708 -72 7375 -10
rect 6881 -81 7044 -72
rect 7212 -81 7375 -72
rect 7428 -224 7486 40
rect 7540 40 7726 96
rect 7772 112 7828 220
rect 7878 158 8052 224
rect 7540 -222 7598 40
rect 7772 36 7950 112
rect 7996 -10 8052 158
rect 8098 40 8164 270
rect 8252 164 8612 222
rect 8270 36 8500 112
rect 8270 -10 8332 36
rect 7665 -72 8332 -10
rect 8556 -23 8612 164
rect 7665 -81 7828 -72
rect 7996 -81 8159 -72
rect 8496 -85 8612 -23
rect 8892 164 9252 222
rect 8892 -23 8948 164
rect 9004 110 9172 112
rect 9004 36 9234 110
rect 9340 40 9406 270
rect 9452 158 9626 224
rect 9172 -10 9234 36
rect 9452 -10 9508 158
rect 9676 112 9732 220
rect 9554 36 9732 112
rect 9778 40 9844 270
rect 10124 40 10190 270
rect 10236 158 10410 224
rect 10236 -10 10292 158
rect 10460 112 10516 220
rect 10338 36 10516 112
rect 10562 40 10628 270
rect 10706 164 11076 222
rect 10734 36 10964 112
rect 10734 -10 10796 36
rect 8892 -85 9008 -23
rect 9172 -72 9839 -10
rect 9345 -81 9508 -72
rect 9676 -81 9839 -72
rect 10129 -72 10796 -10
rect 11020 -23 11076 164
rect 10129 -81 10292 -72
rect 10460 -81 10623 -72
rect 10960 -85 11076 -23
rect 9602 -232 10198 -176
rect 6324 -350 6382 -234
rect 6639 -350 6698 -234
rect 6772 -350 6830 -288
rect 7100 -350 7156 -288
rect 7426 -350 7484 -288
rect 7556 -350 7614 -288
rect 7884 -350 7940 -288
rect 8210 -350 8268 -288
rect 8342 -350 8401 -234
rect 8658 -350 8716 -234
rect 8788 -350 8846 -234
rect 9103 -350 9162 -234
rect 9236 -350 9294 -288
rect 9564 -350 9620 -288
rect 9890 -350 9948 -288
rect 10020 -350 10078 -288
rect 10348 -350 10404 -288
rect 10674 -350 10732 -288
rect 10806 -350 10865 -234
rect 11122 -350 11180 -234
rect 6308 -882 6366 -766
rect 6623 -882 6682 -766
rect 6412 -1032 6528 -1031
rect 6658 -1032 6716 -928
rect 6952 -1026 7018 -914
rect 6412 -1094 6716 -1032
rect 6412 -1280 6468 -1094
rect 6872 -1108 7018 -1026
rect 7234 -976 7864 -930
rect 6872 -1152 6936 -1108
rect 6524 -1228 6936 -1152
rect 7234 -1150 7280 -976
rect 7328 -1072 7400 -1022
rect 6990 -1228 7166 -1154
rect 6412 -1338 6530 -1280
rect 6872 -1296 6936 -1228
rect 7094 -1282 7152 -1228
rect 7234 -1236 7304 -1150
rect 7350 -1252 7400 -1072
rect 7448 -1068 7772 -1022
rect 7448 -1206 7514 -1068
rect 7712 -1084 7772 -1068
rect 7818 -1024 7864 -976
rect 10484 -928 10552 -856
rect 7588 -1252 7654 -1114
rect 7350 -1282 7654 -1252
rect 6308 -1502 6366 -1440
rect 6626 -1502 6684 -1440
rect 6872 -1370 7014 -1296
rect 7094 -1298 7654 -1282
rect 7712 -1286 7766 -1084
rect 7094 -1328 7396 -1298
rect 6948 -1446 7014 -1370
rect 7326 -1446 7396 -1328
rect 7706 -1444 7766 -1286
rect 7818 -1096 8110 -1024
rect 7818 -1286 7864 -1096
rect 8400 -1096 8476 -982
rect 7912 -1240 8194 -1174
rect 8148 -1274 8194 -1240
rect 8428 -1274 8476 -1096
rect 7818 -1332 8098 -1286
rect 8148 -1320 8480 -1274
rect 8030 -1444 8098 -1332
rect 8404 -1438 8480 -1320
rect 9640 -976 10270 -930
rect 9028 -1096 9104 -982
rect 9640 -1024 9686 -976
rect 9028 -1274 9076 -1096
rect 9394 -1096 9686 -1024
rect 9732 -1068 10056 -1022
rect 9732 -1084 9792 -1068
rect 9310 -1240 9592 -1174
rect 9310 -1274 9356 -1240
rect 9024 -1320 9356 -1274
rect 9640 -1286 9686 -1096
rect 9024 -1438 9100 -1320
rect 9406 -1332 9686 -1286
rect 9738 -1286 9792 -1084
rect 9850 -1252 9916 -1114
rect 9990 -1206 10056 -1068
rect 10104 -1072 10176 -1022
rect 10104 -1252 10154 -1072
rect 10224 -1150 10270 -976
rect 10486 -1026 10552 -928
rect 10822 -882 10881 -766
rect 11138 -882 11196 -766
rect 10486 -1108 10632 -1026
rect 10976 -1032 11092 -1031
rect 10778 -1093 11092 -1032
rect 10778 -1094 10985 -1093
rect 10200 -1236 10270 -1150
rect 10568 -1152 10632 -1108
rect 10338 -1228 10514 -1154
rect 10568 -1228 10980 -1152
rect 9850 -1282 10154 -1252
rect 10352 -1282 10410 -1228
rect 9406 -1444 9474 -1332
rect 9738 -1444 9798 -1286
rect 9850 -1298 10410 -1282
rect 10568 -1296 10632 -1228
rect 11036 -1280 11092 -1093
rect 10108 -1328 10410 -1298
rect 10108 -1446 10178 -1328
rect 10490 -1370 10632 -1296
rect 10490 -1446 10556 -1370
rect 10974 -1338 11092 -1280
rect 10820 -1502 10878 -1440
rect 11138 -1502 11196 -1440
<< metal2 >>
rect 6034 2598 6234 2664
rect 6064 1498 6134 2598
rect 7880 2596 8440 2662
rect 8370 2112 8440 2596
rect 8648 2592 8848 2658
rect 8280 1982 8440 2112
rect 8714 1854 8786 2592
rect 9052 2590 9606 2662
rect 11258 2598 11458 2664
rect 9052 2112 9124 2590
rect 9052 1982 9226 2112
rect 7386 1778 10046 1854
rect 7386 1714 7460 1778
rect 9970 1714 10046 1778
rect 7380 1500 7464 1714
rect 9970 1500 10054 1714
rect 6190 -128 6602 -72
rect 6200 -1068 6472 -1012
rect 6196 -1464 6356 -1194
rect 6416 -1300 6472 -1068
rect 6546 -1160 6602 -128
rect 8678 44 8826 922
rect 11358 1666 11430 2598
rect 11352 1498 11430 1666
rect 7912 -1014 9038 -958
rect 7912 -1160 7968 -1014
rect 6546 -1216 7968 -1160
rect 8034 -1216 8386 -1160
rect 8034 -1300 8090 -1216
rect 6416 -1356 8090 -1300
rect 8680 -1464 8828 -1082
rect 8982 -1164 9038 -1014
rect 8982 -1220 9269 -1164
rect 6196 -1614 8828 -1464
<< obsm2 >>
rect 6204 2424 7088 2480
rect 6204 1108 6260 2424
rect 6328 2282 6400 2424
rect 6528 2226 6600 2368
rect 7016 2282 7088 2424
rect 7280 2424 8046 2480
rect 7154 2234 7210 2236
rect 7280 2234 7336 2424
rect 7976 2394 8046 2424
rect 6528 2170 7088 2226
rect 6358 1592 6574 1602
rect 6860 1592 6964 1594
rect 6358 1518 6968 1592
rect 6358 1516 6574 1518
rect 6860 1508 6964 1518
rect 6036 1052 6260 1108
rect 6036 678 6092 1052
rect 7032 932 7088 2170
rect 7154 2178 7336 2234
rect 7496 2226 7568 2368
rect 7976 2282 8048 2394
rect 8176 2226 8248 2368
rect 7154 1040 7210 2178
rect 7496 2170 8248 2226
rect 7496 2106 7568 2170
rect 7266 2050 7568 2106
rect 7266 1184 7322 2050
rect 9450 2424 10326 2480
rect 9250 2226 9320 2368
rect 9450 2282 9520 2424
rect 9934 2226 10004 2368
rect 9250 2170 10214 2226
rect 7630 1592 7740 1600
rect 8018 1592 8220 1604
rect 9282 1592 9476 1604
rect 9766 1592 9874 1600
rect 7630 1518 8234 1592
rect 9270 1518 9874 1592
rect 7630 1516 7740 1518
rect 9766 1516 9874 1518
rect 7266 1128 7430 1184
rect 7154 984 7290 1040
rect 6332 876 7088 932
rect 6332 734 6404 876
rect 6532 678 6604 820
rect 6036 622 6612 678
rect 6556 8 6612 622
rect 6756 562 6812 876
rect 7016 734 7088 876
rect 7234 678 7290 984
rect 7374 932 7430 1128
rect 9014 932 9124 934
rect 10158 932 10214 2170
rect 7374 876 8480 932
rect 7504 678 7576 820
rect 7988 734 8060 876
rect 8192 678 8264 820
rect 7234 622 8328 678
rect 6710 506 6812 562
rect 6710 146 6766 506
rect 8272 142 8328 622
rect 6832 50 7856 106
rect 6832 -184 6888 50
rect 8424 10 8480 876
rect 9014 876 10214 932
rect 9014 354 9070 876
rect 9250 678 9320 820
rect 9450 734 9520 876
rect 9930 678 10000 820
rect 10270 678 10326 2424
rect 10422 2424 11176 2480
rect 10422 2282 10492 2424
rect 10906 2226 10976 2368
rect 10392 2170 10976 2226
rect 11106 2240 11176 2424
rect 11106 2170 11288 2240
rect 10392 932 10448 2170
rect 10556 1592 10660 1594
rect 10928 1592 11114 1602
rect 10544 1518 11114 1592
rect 10556 1508 10660 1518
rect 10928 1516 11114 1518
rect 11232 1074 11288 2170
rect 11232 1024 11292 1074
rect 10390 876 11172 932
rect 10418 734 10488 876
rect 9176 622 10326 678
rect 9014 298 9080 354
rect 9024 4 9080 298
rect 9176 142 9232 622
rect 10676 566 10732 876
rect 10902 678 10972 820
rect 11102 734 11172 876
rect 11236 678 11292 1024
rect 10880 622 11292 678
rect 10676 510 10792 566
rect 9564 268 10406 324
rect 9564 104 9622 268
rect 9566 48 9622 104
rect 6658 -240 6888 -184
rect 6959 -64 7776 -24
rect 9564 -64 9622 48
rect 6959 -80 9622 -64
rect 6658 -1010 6714 -240
rect 6959 -1010 7015 -80
rect 7712 -120 9622 -80
rect 7430 -312 7486 -142
rect 7542 -176 7598 -144
rect 7542 -232 9680 -176
rect 9782 -312 9838 126
rect 10126 -176 10182 126
rect 10348 34 10406 268
rect 10736 138 10792 510
rect 10880 20 10936 622
rect 10114 -232 10544 -176
rect 7430 -368 10408 -312
rect 10352 -1034 10408 -368
rect 10488 -940 10544 -232
rect 10352 -1090 10862 -1034
<< labels >>
rlabel metal2 6064 1498 6134 2598 6 AIN1
port 1 nsew
rlabel metal2 6034 2598 6234 2664 6 AIN1
port 1 nsew
rlabel metal1 6238 872 6284 874 6 AIN1
port 1 nsew
rlabel metal1 6238 874 6292 1258 6 AIN1
port 1 nsew
rlabel metal1 6238 1258 6284 1508 6 AIN1
port 1 nsew
rlabel metal1 6050 1508 6284 1596 6 AIN1
port 1 nsew
rlabel metal1 6238 1596 6284 1862 6 AIN1
port 1 nsew
rlabel metal1 6238 1862 6288 2224 6 AIN1
port 1 nsew
rlabel metal1 6240 2224 6288 2246 6 AIN1
port 1 nsew
rlabel metal1 6064 2578 6134 2580 6 AIN1
port 1 nsew
rlabel metal1 6034 2580 6234 2880 6 AIN1
port 1 nsew
rlabel metal2 8280 1982 8440 2112 6 AIN2
port 2 nsew
rlabel metal2 8370 2112 8440 2596 6 AIN2
port 2 nsew
rlabel metal2 7880 2596 8440 2662 6 AIN2
port 2 nsew
rlabel metal1 8298 868 8344 874 6 AIN2
port 2 nsew
rlabel metal1 8296 874 8344 1258 6 AIN2
port 2 nsew
rlabel metal1 8298 1258 8344 1862 6 AIN2
port 2 nsew
rlabel metal1 8292 1862 8344 1972 6 AIN2
port 2 nsew
rlabel metal1 8292 1972 8358 2124 6 AIN2
port 2 nsew
rlabel metal1 8292 2124 8344 2234 6 AIN2
port 2 nsew
rlabel metal1 8292 2234 8340 2246 6 AIN2
port 2 nsew
rlabel metal1 7908 2576 8108 2878 6 AIN2
port 2 nsew
rlabel metal2 9052 1982 9226 2112 6 AIN3
port 3 nsew
rlabel metal2 9052 2112 9124 2590 6 AIN3
port 3 nsew
rlabel metal2 9052 2590 9606 2662 6 AIN3
port 3 nsew
rlabel metal1 9162 868 9208 874 6 AIN3
port 3 nsew
rlabel metal1 9158 874 9208 1258 6 AIN3
port 3 nsew
rlabel metal1 9162 1258 9208 1862 6 AIN3
port 3 nsew
rlabel metal1 9162 1862 9210 1972 6 AIN3
port 3 nsew
rlabel metal1 9146 1972 9210 2124 6 AIN3
port 3 nsew
rlabel metal1 9162 2124 9210 2246 6 AIN3
port 3 nsew
rlabel metal1 9384 2576 9584 2878 6 AIN3
port 3 nsew
rlabel metal2 11352 1498 11430 1666 6 AIN4
port 4 nsew
rlabel metal2 11358 1666 11430 2598 6 AIN4
port 4 nsew
rlabel metal2 11258 2598 11458 2664 6 AIN4
port 4 nsew
rlabel metal1 11210 874 11258 1258 6 AIN4
port 4 nsew
rlabel metal1 11212 1258 11258 1498 6 AIN4
port 4 nsew
rlabel metal1 11212 1498 11442 1666 6 AIN4
port 4 nsew
rlabel metal1 11212 1666 11258 1862 6 AIN4
port 4 nsew
rlabel metal1 11212 1862 11262 2224 6 AIN4
port 4 nsew
rlabel metal1 11214 2224 11262 2246 6 AIN4
port 4 nsew
rlabel metal1 11258 2578 11458 2880 6 AIN4
port 4 nsew
rlabel metal2 9970 1500 10054 1714 6 AOUT
port 5 nsew
rlabel metal2 7380 1500 7464 1714 6 AOUT
port 5 nsew
rlabel metal2 9970 1714 10046 1778 6 AOUT
port 5 nsew
rlabel metal2 7386 1714 7460 1778 6 AOUT
port 5 nsew
rlabel metal2 7386 1778 10046 1854 6 AOUT
port 5 nsew
rlabel metal2 8714 1854 8786 2592 6 AOUT
port 5 nsew
rlabel metal2 8648 2592 8848 2658 6 AOUT
port 5 nsew
rlabel metal1 10044 868 10090 874 6 AOUT
port 5 nsew
rlabel metal1 7412 868 7458 874 6 AOUT
port 5 nsew
rlabel metal1 10328 874 10376 1258 6 AOUT
port 5 nsew
rlabel metal1 10040 874 10090 1258 6 AOUT
port 5 nsew
rlabel metal1 7412 874 7462 1258 6 AOUT
port 5 nsew
rlabel metal1 7126 874 7174 876 6 AOUT
port 5 nsew
rlabel metal1 10330 1258 10376 1480 6 AOUT
port 5 nsew
rlabel metal1 10044 1258 10090 1480 6 AOUT
port 5 nsew
rlabel metal1 7412 1258 7458 1480 6 AOUT
port 5 nsew
rlabel metal1 7126 876 7180 1258 6 AOUT
port 5 nsew
rlabel metal1 7134 1258 7180 1480 6 AOUT
port 5 nsew
rlabel metal1 9958 1480 10376 1738 6 AOUT
port 5 nsew
rlabel metal1 7134 1480 7476 1738 6 AOUT
port 5 nsew
rlabel metal1 10330 1738 10376 1862 6 AOUT
port 5 nsew
rlabel metal1 10044 1738 10090 1862 6 AOUT
port 5 nsew
rlabel metal1 10330 1862 10380 2238 6 AOUT
port 5 nsew
rlabel metal1 10332 2238 10380 2246 6 AOUT
port 5 nsew
rlabel metal1 10044 1862 10092 2246 6 AOUT
port 5 nsew
rlabel metal1 7412 1738 7458 1862 6 AOUT
port 5 nsew
rlabel metal1 7134 1738 7180 1862 6 AOUT
port 5 nsew
rlabel metal1 7410 1862 7458 2246 6 AOUT
port 5 nsew
rlabel metal1 7122 1862 7180 2238 6 AOUT
port 5 nsew
rlabel metal1 7122 2238 7170 2246 6 AOUT
port 5 nsew
rlabel metal1 8648 2576 8848 2876 6 AOUT
port 5 nsew
rlabel metal2 8982 -1220 9269 -1164 8 SEL[0]
port 6 nsew
rlabel metal2 8982 -1164 9038 -1014 8 SEL[0]
port 6 nsew
rlabel metal2 6546 -1216 7968 -1160 8 SEL[0]
port 6 nsew
rlabel metal2 7912 -1160 7968 -1014 8 SEL[0]
port 6 nsew
rlabel metal2 7912 -1014 9038 -958 8 SEL[0]
port 6 nsew
rlabel metal2 6546 -1160 6602 -128 8 SEL[0]
port 6 nsew
rlabel metal2 6190 -128 6602 -72 8 SEL[0]
port 6 nsew
rlabel metal1 9124 -1228 9258 -1142 8 SEL[0]
port 6 nsew
rlabel metal1 9154 -1142 9258 -1114 8 SEL[0]
port 6 nsew
rlabel metal1 9154 -1114 9348 -1058 8 SEL[0]
port 6 nsew
rlabel metal1 9284 -1058 9348 -978 8 SEL[0]
port 6 nsew
rlabel metal1 9284 -978 9594 -932 8 SEL[0]
port 6 nsew
rlabel metal1 9548 -932 9594 -884 8 SEL[0]
port 6 nsew
rlabel metal1 9548 -884 9644 -838 8 SEL[0]
port 6 nsew
rlabel metal1 5986 -154 6280 -34 8 SEL[0]
port 6 nsew
rlabel metal1 5986 -34 6186 46 6 SEL[0]
port 6 nsew
rlabel metal2 6416 -1356 8090 -1300 8 SEL[1]
port 7 nsew
rlabel metal2 8034 -1300 8090 -1216 8 SEL[1]
port 7 nsew
rlabel metal2 8034 -1216 8386 -1160 8 SEL[1]
port 7 nsew
rlabel metal2 6416 -1300 6472 -1068 8 SEL[1]
port 7 nsew
rlabel metal2 6200 -1068 6472 -1012 8 SEL[1]
port 7 nsew
rlabel metal1 8246 -1228 8380 -1142 8 SEL[1]
port 7 nsew
rlabel metal1 8246 -1142 8350 -1114 8 SEL[1]
port 7 nsew
rlabel metal1 8156 -1114 8350 -1058 8 SEL[1]
port 7 nsew
rlabel metal1 8156 -1058 8220 -978 8 SEL[1]
port 7 nsew
rlabel metal1 5988 -1086 6292 -986 8 SEL[1]
port 7 nsew
rlabel metal1 7910 -978 8220 -932 8 SEL[1]
port 7 nsew
rlabel metal1 7910 -932 7956 -884 8 SEL[1]
port 7 nsew
rlabel metal1 5988 -986 6188 -886 8 SEL[1]
port 7 nsew
rlabel metal1 7860 -884 7956 -838 8 SEL[1]
port 7 nsew
rlabel metal2 6196 -1614 8828 -1464 8 VDD1V8
port 8 nsew
rlabel metal2 8680 -1464 8828 -1082 8 VDD1V8
port 8 nsew
rlabel metal2 6196 -1464 6356 -1194 8 VDD1V8
port 8 nsew
rlabel metal1 8676 -1420 8832 -936 8 VDD1V8
port 8 nsew
rlabel metal1 5982 -1394 6365 -1194 8 VDD1V8
port 8 nsew
rlabel metal1 8266 -936 9238 -886 8 VDD1V8
port 8 nsew
rlabel metal1 8016 -886 9488 -812 8 VDD1V8
port 8 nsew
rlabel metal2 8678 44 8826 922 6 VDD3V3
port 9 nsew
rlabel metal1 10676 -974 10742 -766 8 VDD3V3
port 9 nsew
rlabel metal1 10296 -866 10376 -766 8 VDD3V3
port 9 nsew
rlabel metal1 9922 -884 9988 -766 8 VDD3V3
port 9 nsew
rlabel metal1 7516 -884 7582 -766 8 VDD3V3
port 9 nsew
rlabel metal1 7128 -866 7208 -766 8 VDD3V3
port 9 nsew
rlabel metal1 6762 -974 6828 -766 8 VDD3V3
port 9 nsew
rlabel metal1 6272 -766 11232 -606 8 VDD3V3
port 9 nsew
rlabel metal1 10760 -606 10976 -510 8 VDD3V3
port 9 nsew
rlabel metal1 8678 -606 8826 -510 8 VDD3V3
port 9 nsew
rlabel metal1 6528 -606 6744 -510 8 VDD3V3
port 9 nsew
rlabel metal1 6288 -510 11216 -350 8 VDD3V3
port 9 nsew
rlabel metal1 8716 -350 8788 -234 8 VDD3V3
port 9 nsew
rlabel metal1 8678 -234 8826 226 8 VDD3V3
port 9 nsew
rlabel metal1 8976 1794 9052 1840 6 VDD3V3
port 9 nsew
rlabel metal1 11358 1840 11406 1852 6 VDD3V3
port 9 nsew
rlabel metal1 11358 1852 11468 2424 6 VDD3V3
port 9 nsew
rlabel metal1 10674 1840 10722 1842 6 VDD3V3
port 9 nsew
rlabel metal1 10188 1840 10236 1842 6 VDD3V3
port 9 nsew
rlabel metal1 10672 1842 10722 2268 6 VDD3V3
port 9 nsew
rlabel metal1 10186 1842 10236 2268 6 VDD3V3
port 9 nsew
rlabel metal1 9702 1840 9750 1844 6 VDD3V3
port 9 nsew
rlabel metal1 9690 1844 9750 2268 6 VDD3V3
port 9 nsew
rlabel metal1 8976 1840 9066 2268 6 VDD3V3
port 9 nsew
rlabel metal1 10672 2268 10718 2424 6 VDD3V3
port 9 nsew
rlabel metal1 10186 2268 10232 2424 6 VDD3V3
port 9 nsew
rlabel metal1 9690 2268 9736 2424 6 VDD3V3
port 9 nsew
rlabel metal1 8976 2268 9052 2424 6 VDD3V3
port 9 nsew
rlabel metal1 8680 786 8822 2424 6 VDD3V3
port 9 nsew
rlabel metal1 8436 1794 8514 2424 6 VDD3V3
port 9 nsew
rlabel metal1 7752 1840 7800 1844 6 VDD3V3
port 9 nsew
rlabel metal1 7752 1844 7806 2268 6 VDD3V3
port 9 nsew
rlabel metal1 7266 1840 7314 1842 6 VDD3V3
port 9 nsew
rlabel metal1 7260 1842 7314 2268 6 VDD3V3
port 9 nsew
rlabel metal1 6780 1840 6828 2268 6 VDD3V3
port 9 nsew
rlabel metal1 6096 1840 6144 1846 6 VDD3V3
port 9 nsew
rlabel metal1 6094 1846 6144 2268 6 VDD3V3
port 9 nsew
rlabel metal1 7760 2268 7806 2424 6 VDD3V3
port 9 nsew
rlabel metal1 7260 2268 7306 2424 6 VDD3V3
port 9 nsew
rlabel metal1 6780 2268 6826 2424 6 VDD3V3
port 9 nsew
rlabel metal1 6094 2268 6140 2424 6 VDD3V3
port 9 nsew
rlabel metal1 6094 2424 11468 2530 6 VDD3V3
port 9 nsew
rlabel metal1 7174 2530 7374 2870 6 VDD3V3
port 9 nsew
rlabel metal1 11304 -1664 11464 -1662 8 VSSA
port 10 nsew
rlabel metal1 6272 -1662 11464 -1502 8 VSSA
port 10 nsew
rlabel metal1 11304 -1502 11464 590 8 VSSA
port 10 nsew
rlabel metal1 10680 -1502 10744 -1326 8 VSSA
port 10 nsew
rlabel metal1 10300 -1502 10370 -1374 8 VSSA
port 10 nsew
rlabel metal1 9920 -1502 9990 -1344 8 VSSA
port 10 nsew
rlabel metal1 9536 -1502 9622 -1382 8 VSSA
port 10 nsew
rlabel metal1 9218 -1502 9282 -1366 8 VSSA
port 10 nsew
rlabel metal1 8222 -1502 8286 -1366 8 VSSA
port 10 nsew
rlabel metal1 7882 -1502 7968 -1382 8 VSSA
port 10 nsew
rlabel metal1 7514 -1502 7584 -1344 8 VSSA
port 10 nsew
rlabel metal1 7134 -1502 7204 -1374 8 VSSA
port 10 nsew
rlabel metal1 6760 -1502 6824 -1326 8 VSSA
port 10 nsew
rlabel metal1 5994 384 6324 386 6 VSSA
port 10 nsew
rlabel metal1 5994 386 11216 546 6 VSSA
port 10 nsew
rlabel metal1 10962 546 11216 590 6 VSSA
port 10 nsew
rlabel metal1 10962 590 11464 592 6 VSSA
port 10 nsew
rlabel metal1 9330 546 9494 592 6 VSSA
port 10 nsew
rlabel metal1 7998 546 8164 592 6 VSSA
port 10 nsew
rlabel metal1 5994 546 6516 592 6 VSSA
port 10 nsew
rlabel metal1 5994 592 11464 696 6 VSSA
port 10 nsew
rlabel metal1 11358 696 11464 852 6 VSSA
port 10 nsew
rlabel metal1 10676 696 10722 852 6 VSSA
port 10 nsew
rlabel metal1 10194 696 10240 852 6 VSSA
port 10 nsew
rlabel metal1 9698 696 9744 852 6 VSSA
port 10 nsew
rlabel metal1 11354 852 11464 1266 6 VSSA
port 10 nsew
rlabel metal1 11354 1266 11402 1280 6 VSSA
port 10 nsew
rlabel metal1 10820 864 10866 874 6 VSSA
port 10 nsew
rlabel metal1 10814 874 10866 978 6 VSSA
port 10 nsew
rlabel metal1 10670 852 10722 978 6 VSSA
port 10 nsew
rlabel metal1 10670 978 10866 1094 6 VSSA
port 10 nsew
rlabel metal1 10814 1094 10866 1258 6 VSSA
port 10 nsew
rlabel metal1 10820 1258 10866 1862 6 VSSA
port 10 nsew
rlabel metal1 10670 1094 10722 1270 6 VSSA
port 10 nsew
rlabel metal1 10184 852 10240 1260 6 VSSA
port 10 nsew
rlabel metal1 10670 1270 10718 1280 6 VSSA
port 10 nsew
rlabel metal1 10184 1260 10232 1280 6 VSSA
port 10 nsew
rlabel metal1 9698 852 9746 1024 6 VSSA
port 10 nsew
rlabel metal1 9016 696 9062 852 6 VSSA
port 10 nsew
rlabel metal1 8444 696 8490 852 6 VSSA
port 10 nsew
rlabel metal1 7752 696 7798 852 6 VSSA
port 10 nsew
rlabel metal1 7270 696 7316 852 6 VSSA
port 10 nsew
rlabel metal1 6776 696 6822 852 6 VSSA
port 10 nsew
rlabel metal1 6092 696 6146 852 6 VSSA
port 10 nsew
rlabel metal1 9556 870 9602 874 6 VSSA
port 10 nsew
rlabel metal1 9554 874 9602 1024 6 VSSA
port 10 nsew
rlabel metal1 9554 1024 9746 1122 6 VSSA
port 10 nsew
rlabel metal1 9698 1122 9746 1280 6 VSSA
port 10 nsew
rlabel metal1 9554 1122 9602 1258 6 VSSA
port 10 nsew
rlabel metal1 9556 1258 9602 1862 6 VSSA
port 10 nsew
rlabel metal1 9014 852 9062 1280 6 VSSA
port 10 nsew
rlabel metal1 8440 852 8490 1264 6 VSSA
port 10 nsew
rlabel metal1 7896 870 7942 874 6 VSSA
port 10 nsew
rlabel metal1 7896 874 7948 1024 6 VSSA
port 10 nsew
rlabel metal1 7752 852 7804 1024 6 VSSA
port 10 nsew
rlabel metal1 7752 1024 7948 1122 6 VSSA
port 10 nsew
rlabel metal1 7896 1122 7948 1258 6 VSSA
port 10 nsew
rlabel metal1 8440 1264 8488 1280 6 VSSA
port 10 nsew
rlabel metal1 7896 1258 7942 1862 6 VSSA
port 10 nsew
rlabel metal1 7752 1122 7804 1266 6 VSSA
port 10 nsew
rlabel metal1 7756 1266 7804 1280 6 VSSA
port 10 nsew
rlabel metal1 7270 852 7318 1280 6 VSSA
port 10 nsew
rlabel metal1 6776 852 6832 978 6 VSSA
port 10 nsew
rlabel metal1 6640 864 6686 874 6 VSSA
port 10 nsew
rlabel metal1 6640 874 6688 978 6 VSSA
port 10 nsew
rlabel metal1 6640 978 6832 1094 6 VSSA
port 10 nsew
rlabel metal1 6776 1094 6832 1270 6 VSSA
port 10 nsew
rlabel metal1 6640 1094 6688 1258 6 VSSA
port 10 nsew
rlabel metal1 6784 1270 6832 1280 6 VSSA
port 10 nsew
rlabel metal1 10818 1862 10866 2246 6 VSSA
port 10 nsew
rlabel metal1 9556 1862 9606 2234 6 VSSA
port 10 nsew
rlabel metal1 9558 2234 9606 2246 6 VSSA
port 10 nsew
rlabel metal1 7896 1862 7944 2246 6 VSSA
port 10 nsew
rlabel metal1 6640 1258 6686 1862 6 VSSA
port 10 nsew
rlabel metal1 6092 852 6148 1278 6 VSSA
port 10 nsew
rlabel metal1 6100 1278 6148 1280 6 VSSA
port 10 nsew
rlabel metal1 6636 1862 6686 2230 6 VSSA
port 10 nsew
rlabel metal1 6636 2230 6684 2246 6 VSSA
port 10 nsew
<< properties >>
string LEFview TRUE
string FIXED_BBOX 5982 -1710 11512 2880
string GDS_FILE ~/design/ip/AMUX4_3V/11.0/gds/AMUX4_3V.gds
string GDS_START 28490
string GDS_END 58642
<< end >>
