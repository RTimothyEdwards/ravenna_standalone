magic
tech EFXH018D
magscale 1 2
timestamp 1569591303
<< error_s >>
rect 32100 406800 32500 413600
rect 48900 406800 49300 413600
rect 65700 406800 66100 413600
rect 82500 406800 82900 413600
rect 99300 406800 99700 413600
rect 116100 406800 116500 413600
rect 132900 406800 133300 413600
rect 149700 406800 150100 413600
rect 159700 406800 160100 413600
rect 169700 406800 170100 413600
rect 179700 406800 180100 413600
rect 189700 406800 190100 413600
rect 206500 406800 206900 413600
rect 223300 406800 223700 413600
rect 233300 406800 233700 413600
rect 250100 406800 250500 413600
rect 266900 406800 267300 413600
rect 283700 406800 284100 413600
rect 293700 406800 294100 413600
rect 303700 406800 304100 413600
rect 313700 406800 314100 413600
rect 323700 406800 324100 413600
rect 333500 406800 334200 413600
rect 333792 406708 334200 406800
rect 333600 406300 334200 406708
rect 425600 406708 426008 413600
rect 426100 406800 426700 413600
rect 443100 406800 443500 413600
rect 459900 406800 460300 413600
rect 463900 406800 464300 413600
rect 465900 406800 466300 413600
rect 482700 406800 483100 413600
rect 425600 406300 426200 406708
rect 344122 402287 349406 402695
rect 344122 395944 344530 402287
rect 344622 401787 348906 402195
rect 344622 396444 345030 401787
rect 345435 396633 347730 401225
rect 348498 396444 348906 401787
rect 344622 396036 348906 396444
rect 348998 395944 349406 402287
rect 344122 395536 349406 395944
rect 410394 402019 415544 402427
rect 410394 395944 410802 402019
rect 410894 401519 415044 401927
rect 410894 396444 411302 401519
rect 411805 396633 414100 401225
rect 414636 396444 415044 401519
rect 410894 396036 415044 396444
rect 415136 395944 415544 402019
rect 410394 395536 415544 395944
rect 429176 392456 429180 405896
rect 445976 392456 445980 405896
rect 35048 392440 45704 392456
rect 51848 392440 62504 392456
rect 68648 392440 79304 392456
rect 85448 392440 96000 392456
rect 102248 392440 112904 392456
rect 119048 392440 129704 392456
rect 135848 392440 146504 392456
rect 192632 392440 203288 392456
rect 209432 392440 220088 392456
rect 236312 392440 246968 392456
rect 253112 392440 263768 392456
rect 269800 392440 280456 392456
rect 429176 392440 439944 392456
rect 445976 392440 456744 392456
rect 333600 391668 334200 392076
rect 333792 391576 334200 391668
rect 32100 385176 32500 391576
rect 48900 385176 49300 391576
rect 65700 385176 66100 391576
rect 82500 385176 82900 391576
rect 99300 385176 99700 391576
rect 116100 385176 116500 391576
rect 132900 385176 133300 391576
rect 149700 385176 150100 391576
rect 159700 385176 160100 391576
rect 169700 385176 170100 391576
rect 179700 385176 180100 391576
rect 189700 385176 190100 391576
rect 206500 385176 206900 391576
rect 223300 385176 223700 391576
rect 233300 385176 233700 391576
rect 250100 385176 250500 391576
rect 266900 385176 267300 391576
rect 283700 385176 284100 391576
rect 293700 385176 294100 391576
rect 303700 385176 304100 391576
rect 313700 385176 314100 391576
rect 323700 385176 324100 391576
rect 333500 385235 334200 391576
rect 333000 385176 334200 385235
rect 333000 385084 333700 385176
rect 333792 385084 334200 385176
rect 333000 384923 334200 385084
rect 333000 384831 333700 384923
rect 333792 384831 334200 384923
rect 31900 383948 32500 384676
rect 48700 383948 49300 384676
rect 65500 383948 66100 384676
rect 82300 383948 82900 384676
rect 99100 383948 99700 384676
rect 115900 383948 116500 384676
rect 132700 383948 133300 384676
rect 149500 383948 150100 384676
rect 159500 383948 160100 384676
rect 169500 383948 170100 384676
rect 179500 383948 180100 384676
rect 189500 383948 190100 384676
rect 206300 383948 206900 384676
rect 223100 383948 223700 384676
rect 233100 383948 233700 384676
rect 249900 383948 250500 384676
rect 266700 383948 267300 384676
rect 283500 383948 284100 384676
rect 293500 383948 294100 384676
rect 303500 383948 304100 384676
rect 313500 383948 314100 384676
rect 323500 383948 324100 384676
rect 333000 384359 334200 384831
rect 333500 383948 334200 384359
rect 333600 383667 334200 383948
rect 333000 383587 334200 383667
rect 333000 383467 333700 383587
rect 333792 383467 334200 383587
rect 31900 382848 32500 383448
rect 48700 382848 49300 383448
rect 65500 382848 66100 383448
rect 82300 382848 82900 383448
rect 99100 382848 99700 383448
rect 115900 382848 116500 383448
rect 132700 382848 133300 383448
rect 149500 382848 150100 383448
rect 159500 382848 160100 383448
rect 169500 382848 170100 383448
rect 179500 382848 180100 383448
rect 189500 382848 190100 383448
rect 206300 382848 206900 383448
rect 223100 382848 223700 383448
rect 233100 382848 233700 383448
rect 249900 382848 250500 383448
rect 266700 382848 267300 383448
rect 283500 382848 284100 383448
rect 293500 382848 294100 383448
rect 303500 382848 304100 383448
rect 313500 382848 314100 383448
rect 323500 382848 324100 383448
rect 333000 383067 334200 383467
rect 333500 382848 334200 383067
rect 333600 382547 334200 382848
rect 333792 382428 334200 382547
rect 333600 382348 334200 382428
rect 0 381700 6800 382100
rect 22024 381700 28424 382100
rect 28924 381500 29652 382100
rect 30152 381500 30752 382100
rect 31252 381500 31852 382100
rect 31900 381748 32500 382348
rect 48700 381748 49300 382348
rect 65500 381748 66100 382348
rect 82300 381748 82900 382348
rect 99100 381748 99700 382348
rect 115900 381748 116500 382348
rect 132700 381748 133300 382348
rect 149500 381748 150100 382348
rect 159500 381748 160100 382348
rect 169500 381748 170100 382348
rect 179500 381748 180100 382348
rect 189500 381748 190100 382348
rect 206300 381748 206900 382348
rect 223100 381748 223700 382348
rect 233100 381748 233700 382348
rect 249900 381748 250500 382348
rect 266700 381748 267300 382348
rect 283500 381748 284100 382348
rect 293500 381748 294100 382348
rect 303500 381748 304100 382348
rect 313500 381748 314100 382348
rect 323500 381748 324100 382348
rect 333500 381748 334200 382348
rect 333792 381656 334200 381748
rect 333600 381443 334200 381656
rect 425600 391668 426200 392076
rect 425600 385084 426008 391668
rect 426100 385235 426700 391576
rect 426100 385084 426800 385235
rect 443100 385176 443500 391576
rect 459900 385176 460300 391576
rect 463900 385176 464300 391576
rect 465900 385176 466300 391576
rect 482700 385176 483100 391576
rect 425600 384923 426800 385084
rect 425600 384548 426008 384923
rect 426100 384548 426800 384923
rect 425600 384267 426800 384548
rect 425600 383948 426700 384267
rect 442900 383948 443500 384676
rect 459700 383948 460300 384676
rect 463700 383948 464300 384676
rect 465700 383948 466300 384676
rect 482500 383948 483100 384676
rect 425600 383448 426008 383948
rect 426100 383667 426700 383948
rect 426100 383448 426800 383667
rect 425600 382947 426800 383448
rect 425600 382848 426700 382947
rect 442900 382848 443500 383448
rect 459700 382848 460300 383448
rect 463700 382848 464300 383448
rect 465700 382848 466300 383448
rect 482500 382848 483100 383448
rect 425600 381656 426008 382848
rect 426100 382547 426700 382848
rect 426100 381748 426700 382428
rect 442900 381748 443500 382348
rect 459700 381748 460300 382348
rect 463700 381748 464300 382348
rect 465700 381748 466300 382348
rect 482500 382100 483100 382348
rect 482500 381748 483348 382100
rect 425600 381443 426200 381656
rect 482748 381500 483348 381748
rect 483848 381500 484448 382100
rect 484948 381500 485676 382100
rect 486176 381700 492576 382100
rect 507800 381700 514600 382100
rect 0 364900 6800 365300
rect 22024 364900 28424 365300
rect 28924 364700 29652 365300
rect 30152 364700 30752 365300
rect 31252 364700 31852 365300
rect 482748 364700 483348 365300
rect 483848 364700 484448 365300
rect 484948 364700 485676 365300
rect 486176 364900 492576 365300
rect 507800 364900 514600 365300
rect 334216 363026 340056 363100
rect 334216 362980 334290 363026
rect 339982 362920 340056 363026
rect 340428 363026 346268 363100
rect 340428 362980 340502 363026
rect 346194 362920 346268 363026
rect 0 348100 6800 348500
rect 22024 348100 28424 348500
rect 28924 347900 29652 348500
rect 30152 347900 30752 348500
rect 31252 347900 31852 348500
rect 482748 347900 483348 348500
rect 483848 347900 484448 348500
rect 484948 347900 485676 348500
rect 486176 348100 492576 348500
rect 507800 348100 514600 348500
rect 0 338100 6800 338500
rect 22024 338100 28424 338500
rect 28924 337900 29652 338500
rect 30152 337900 30752 338500
rect 31252 337900 31852 338500
rect 482748 331100 483348 331700
rect 483848 331100 484448 331700
rect 484948 331100 485676 331700
rect 486176 331300 492576 331700
rect 507800 331300 514600 331700
rect 0 321300 6800 321700
rect 22024 321300 28424 321700
rect 28924 321100 29652 321700
rect 30152 321100 30752 321700
rect 31252 321100 31852 321700
rect 482748 314300 483348 314900
rect 483848 314300 484448 314900
rect 484948 314300 485676 314900
rect 486176 314500 492576 314900
rect 507800 314500 514600 314900
rect 62854 312560 62922 312679
rect 63186 312560 63244 312678
rect 0 304500 6800 304900
rect 22024 304500 28424 304900
rect 28924 304300 29652 304900
rect 30152 304300 30752 304900
rect 31252 304300 31852 304900
rect 482748 297500 483348 298100
rect 483848 297500 484448 298100
rect 484948 297500 485676 298100
rect 486176 297700 492576 298100
rect 507800 297700 514600 298100
rect 0 287700 6800 288100
rect 22024 287700 28424 288100
rect 28924 287500 29652 288100
rect 30152 287500 30752 288100
rect 31252 287500 31852 288100
rect 482748 287500 483348 288100
rect 483848 287500 484448 288100
rect 484948 287500 485676 288100
rect 486176 287700 492576 288100
rect 507800 287700 514600 288100
rect 482748 277500 483348 278100
rect 483848 277500 484448 278100
rect 484948 277500 485676 278100
rect 486176 277700 492576 278100
rect 507800 277700 514600 278100
rect 7720 273720 21064 273780
rect 0 270900 6800 271300
rect 22024 270900 28424 271300
rect 28924 270700 29652 271300
rect 30152 270700 30752 271300
rect 31252 270700 31852 271300
rect 482748 267500 483348 268100
rect 483848 267500 484448 268100
rect 484948 267500 485676 268100
rect 486176 267700 492576 268100
rect 507800 267700 514600 268100
rect 30152 260300 30752 260900
rect 31252 260300 31852 260900
rect 0 258500 6800 258900
rect 22024 258500 28424 258900
rect 28924 258300 29652 258900
rect 30152 258300 30752 258900
rect 31252 258300 31852 258900
rect 482748 257500 483348 258100
rect 483848 257500 484448 258100
rect 484948 257500 485676 258100
rect 486176 257700 492576 258100
rect 507800 257700 514600 258100
rect 0 241700 6800 242100
rect 22024 241700 28424 242100
rect 28924 241500 29652 242100
rect 30152 241500 30752 242100
rect 31252 241500 31852 242100
rect 482748 240700 483348 241300
rect 483848 240700 484448 241300
rect 484948 240700 485676 241300
rect 486176 240900 492576 241300
rect 507800 240900 514600 241300
rect 0 224900 6800 225300
rect 22024 224900 28424 225300
rect 28924 224700 29652 225300
rect 30152 224700 30752 225300
rect 31252 224700 31852 225300
rect 482748 223900 483348 224500
rect 483848 223900 484448 224500
rect 484948 223900 485676 224500
rect 486176 224100 492576 224500
rect 507800 224100 514600 224500
rect 482748 213900 483348 214500
rect 483848 213900 484448 214500
rect 484948 213900 485676 214500
rect 486176 214100 492576 214500
rect 507800 214100 514600 214500
rect 0 208100 6800 208500
rect 22024 208100 28424 208500
rect 28924 207900 29652 208500
rect 30152 207900 30752 208500
rect 31252 207900 31852 208500
rect 482748 197100 483348 197700
rect 483848 197100 484448 197700
rect 484948 197100 485676 197700
rect 486176 197300 492576 197700
rect 507800 197300 514600 197700
rect 0 191300 6800 191700
rect 22024 191300 28424 191700
rect 28924 191100 29652 191700
rect 30152 191100 30752 191700
rect 31252 191100 31852 191700
rect 482748 180300 483348 180900
rect 483848 180300 484448 180900
rect 484948 180300 485676 180900
rect 486176 180500 492576 180900
rect 507800 180500 514600 180900
rect 0 174500 6800 174900
rect 22024 174500 28424 174900
rect 28924 174300 29652 174900
rect 30152 174300 30752 174900
rect 31252 174300 31852 174900
rect 482748 170300 483348 170900
rect 483848 170300 484448 170900
rect 484948 170300 485676 170900
rect 486176 170500 492576 170900
rect 507800 170500 514600 170900
rect 482748 160300 483348 160900
rect 483848 160300 484448 160900
rect 484948 160300 485676 160900
rect 486176 160500 492576 160900
rect 507800 160500 514600 160900
rect 0 157700 6800 158100
rect 22024 157700 28424 158100
rect 28924 157500 29652 158100
rect 30152 157500 30752 158100
rect 31252 157500 31852 158100
rect 482748 150300 483348 150900
rect 483848 150300 484448 150900
rect 484948 150300 485676 150900
rect 486176 150500 492576 150900
rect 507800 150500 514600 150900
rect 0 140900 6800 141300
rect 22024 140900 28424 141300
rect 28924 140700 29652 141300
rect 30152 140700 30752 141300
rect 31252 140700 31852 141300
rect 482748 133500 483348 134100
rect 483848 133500 484448 134100
rect 484948 133500 485676 134100
rect 486176 133700 492576 134100
rect 507800 133700 514600 134100
rect 0 130900 6800 131300
rect 22024 130900 28424 131300
rect 28924 130700 29652 131300
rect 30152 130700 30752 131300
rect 31252 130700 31852 131300
rect 482748 116700 483348 117300
rect 483848 116700 484448 117300
rect 484948 116700 485676 117300
rect 486176 116900 492576 117300
rect 507800 116900 514600 117300
rect 28365 114400 31253 114600
rect 0 113800 6800 114400
rect 22024 114000 31852 114400
rect 6892 113708 7300 114000
rect 0 113300 7300 113708
rect 21524 113708 21932 114000
rect 22024 113800 28424 114000
rect 28516 113708 28677 114000
rect 28769 113800 30013 114000
rect 30133 113800 31852 114000
rect 21524 113300 31882 113708
rect 63396 109056 63464 109064
rect 63684 109056 63752 109064
rect 63972 109056 64040 109064
rect 64260 109056 64263 109064
rect 61662 108231 61730 108347
rect 62018 108231 62076 108293
rect 12191 107332 16828 107740
rect 12191 104048 12599 107332
rect 12691 106832 16328 107240
rect 12691 104548 13099 106832
rect 15920 104548 16328 106832
rect 12691 104140 16328 104548
rect 16420 104048 16828 107332
rect 482748 106700 483348 107300
rect 483848 106700 484448 107300
rect 484948 106700 485676 107300
rect 486176 106900 492576 107300
rect 507800 106900 514600 107300
rect 12191 103640 16828 104048
rect 482748 96700 483348 97300
rect 483848 96700 484448 97300
rect 484948 96700 485676 97300
rect 486176 96900 492576 97300
rect 507800 96900 514600 97300
rect 482748 86700 483348 87300
rect 483848 86700 484448 87300
rect 484948 86700 485676 87300
rect 486176 86900 492576 87300
rect 507800 86900 514600 87300
rect 482748 76700 483348 77300
rect 483848 76700 484448 77300
rect 484948 76700 485676 77300
rect 486176 76900 492576 77300
rect 507800 76900 514600 77300
rect 11773 68692 17007 69100
rect 11773 65168 12181 68692
rect 12273 68192 16507 68600
rect 12273 65668 12681 68192
rect 16099 65668 16507 68192
rect 12273 65260 16507 65668
rect 16599 65168 17007 68692
rect 11773 64760 17007 65168
rect 482748 59900 483348 60500
rect 483848 59900 484448 60500
rect 484948 59900 485676 60500
rect 486176 60100 492576 60500
rect 507800 60100 514600 60500
rect 0 59092 7300 59500
rect 0 58700 6800 59092
rect 6892 58800 7300 59092
rect 21524 59092 31882 59500
rect 21524 58800 21932 59092
rect 22024 58700 28424 59092
rect 28516 58800 28677 59092
rect 28769 58800 30013 59092
rect 30133 59000 31053 59092
rect 31172 59000 31852 59092
rect 30133 58800 31852 59000
rect 28924 58700 29652 58800
rect 30152 58700 30752 58800
rect 31252 58700 31852 58800
rect 198932 50574 199006 50680
rect 204698 50574 204772 50620
rect 198932 50500 204772 50574
rect 205144 50574 205218 50620
rect 210910 50574 210984 50680
rect 205144 50500 210984 50574
rect 482748 43100 483348 43700
rect 483848 43100 484448 43700
rect 484948 43100 485676 43700
rect 486176 43300 492576 43700
rect 507800 43300 514600 43700
rect 0 42100 6800 42500
rect 22024 42100 28424 42500
rect 28924 41900 29652 42500
rect 30152 41900 30752 42500
rect 31252 41900 31852 42500
rect 482748 32900 483348 33500
rect 483848 32900 484448 33500
rect 484948 32900 485676 33500
rect 486176 33300 492576 33500
rect 507800 33300 514600 33500
rect 0 32100 6800 32500
rect 22024 32100 28424 32500
rect 28924 31900 29652 32500
rect 30152 31900 30752 32500
rect 31252 31900 31852 32500
rect 119000 31944 119600 32157
rect 119192 31852 119600 31944
rect 31900 31252 32500 31852
rect 32900 31252 33500 31852
rect 34000 31252 34600 31852
rect 50700 31252 51300 31852
rect 67500 31252 68100 31852
rect 84300 31252 84900 31852
rect 101100 31252 101700 31852
rect 117900 31252 118500 31852
rect 119000 31172 119600 31852
rect 119000 31053 119100 31172
rect 119192 31053 119600 31172
rect 31900 30152 32500 30752
rect 32900 30152 33500 30752
rect 34000 30152 34600 30752
rect 50700 30152 51300 30752
rect 67500 30152 68100 30752
rect 84300 30152 84900 30752
rect 101100 30152 101700 30752
rect 117900 30152 118500 30752
rect 119000 30653 119600 31053
rect 119000 30533 119100 30653
rect 119192 30533 119600 30653
rect 119000 30133 119600 30533
rect 119192 30013 119600 30133
rect 31900 28924 32500 29652
rect 32900 28924 33500 29652
rect 34000 28924 34600 29652
rect 50700 28924 51300 29652
rect 67500 28924 68100 29652
rect 84300 28924 84900 29652
rect 101100 28924 101700 29652
rect 117900 28924 118500 29652
rect 119000 29333 119600 30013
rect 119000 29241 119100 29333
rect 119192 29241 119600 29333
rect 119000 29057 119600 29241
rect 119000 28965 119100 29057
rect 119192 28965 119600 29057
rect 119000 28769 119600 28965
rect 119192 28677 119600 28769
rect 119000 28516 119600 28677
rect 119192 28424 119600 28516
rect 32100 22024 32500 28424
rect 33000 22024 33500 28424
rect 34100 22024 34600 28424
rect 50900 22024 51300 28424
rect 67700 22024 68100 28424
rect 84500 22024 84900 28424
rect 101300 22024 101700 28424
rect 118000 22024 118500 28424
rect 119000 22024 119600 28424
rect 119192 21932 119600 22024
rect 119000 21524 119600 21932
rect 211000 31944 211600 32157
rect 211000 31852 211408 31944
rect 482748 31900 483348 32500
rect 483848 31900 484448 32500
rect 484948 31900 485676 32500
rect 486176 32100 492576 32500
rect 507800 32100 514600 32500
rect 211000 31252 212100 31852
rect 219500 31252 220100 31852
rect 220500 31252 221100 31852
rect 230500 31252 231100 31852
rect 247300 31252 247900 31852
rect 257300 31252 257900 31852
rect 267300 31252 267900 31852
rect 284100 31252 284700 31852
rect 300900 31252 301500 31852
rect 310900 31252 311500 31852
rect 327700 31252 328300 31852
rect 344500 31252 345100 31852
rect 354500 31252 355100 31852
rect 364500 31252 365100 31852
rect 381300 31252 381900 31852
rect 398100 31252 398700 31852
rect 414900 31252 415500 31852
rect 431700 31252 432300 31852
rect 448500 31252 449100 31852
rect 458500 31252 459100 31852
rect 462500 31252 463100 31852
rect 464500 31252 465100 31852
rect 465500 31252 466100 31852
rect 482500 31252 483100 31852
rect 211000 30752 211408 31252
rect 211500 30752 212200 31252
rect 211000 30533 212200 30752
rect 211000 30152 212100 30533
rect 219500 30152 220100 30752
rect 220500 30152 221100 30752
rect 230500 30152 231100 30752
rect 247300 30152 247900 30752
rect 257300 30152 257900 30752
rect 267300 30152 267900 30752
rect 284100 30152 284700 30752
rect 300900 30152 301500 30752
rect 310900 30152 311500 30752
rect 327700 30152 328300 30752
rect 344500 30152 345100 30752
rect 354500 30152 355100 30752
rect 364500 30152 365100 30752
rect 381300 30152 381900 30752
rect 398100 30152 398700 30752
rect 414900 30152 415500 30752
rect 431700 30152 432300 30752
rect 448500 30152 449100 30752
rect 458500 30152 459100 30752
rect 462500 30152 463100 30752
rect 464500 30152 465100 30752
rect 465500 30152 466100 30752
rect 482500 30152 483100 30752
rect 211000 29524 211408 30152
rect 211500 30133 212100 30152
rect 211500 29933 212100 30013
rect 211500 29524 212200 29933
rect 211000 28965 212200 29524
rect 211000 28924 212100 28965
rect 219500 28924 220100 29652
rect 220500 28924 221100 29652
rect 230500 28924 231100 29652
rect 247300 28924 247900 29652
rect 257300 28924 257900 29652
rect 267300 28924 267900 29652
rect 284100 28924 284700 29652
rect 300900 28924 301500 29652
rect 310900 28924 311500 29652
rect 327700 28924 328300 29652
rect 344500 28924 345100 29652
rect 354500 28924 355100 29652
rect 364500 28924 365100 29652
rect 381300 28924 381900 29652
rect 398100 28924 398700 29652
rect 414900 28924 415500 29652
rect 431700 28924 432300 29652
rect 448500 28924 449100 29652
rect 458500 28924 459100 29652
rect 462500 28924 463100 29652
rect 464500 28924 465100 29652
rect 465500 28924 466100 29652
rect 482500 28924 483100 29652
rect 211000 28677 211408 28924
rect 211500 28769 212100 28924
rect 211000 28516 211600 28677
rect 211000 21932 211408 28516
rect 211500 22024 212100 28424
rect 219700 22024 220100 28424
rect 220700 22024 221100 28424
rect 230700 22024 231100 28424
rect 247500 22024 247900 28424
rect 257500 22024 257900 28424
rect 267500 22024 267900 28424
rect 284300 22024 284700 28424
rect 301100 22024 301500 28424
rect 311100 22024 311500 28424
rect 327900 22024 328300 28424
rect 344700 22024 345100 28424
rect 354700 22024 355100 28424
rect 364700 22024 365100 28424
rect 381500 22024 381900 28424
rect 398300 22024 398700 28424
rect 415100 22024 415500 28424
rect 431900 22024 432300 28424
rect 448700 22024 449100 28424
rect 458700 22024 459100 28424
rect 462700 22024 463100 28424
rect 464700 22024 465100 28424
rect 465900 22024 466100 28424
rect 482700 22024 483100 28424
rect 211000 21524 211600 21932
rect 129656 17656 134806 18064
rect 129656 11581 130064 17656
rect 130156 17156 134306 17564
rect 130156 12081 130564 17156
rect 130818 12162 133191 16645
rect 133898 12081 134306 17156
rect 130156 11673 134306 12081
rect 134398 11581 134806 17656
rect 129656 11173 134806 11581
rect 195794 17656 201078 18064
rect 195794 11313 196202 17656
rect 196294 17156 200578 17564
rect 196294 11813 196702 17156
rect 197145 12162 199650 16777
rect 200170 11813 200578 17156
rect 196294 11405 200578 11813
rect 200670 11313 201078 17656
rect 195794 10905 201078 11313
rect 287160 7720 287180 21064
rect 367576 7720 367580 21064
rect 384376 7720 384380 21064
rect 401176 7720 401180 21064
rect 417976 7720 417980 21064
rect 119000 6892 119600 7300
rect 119192 6800 119600 6892
rect 32100 0 32500 6800
rect 33000 0 33500 6800
rect 34100 0 34600 6800
rect 50900 0 51300 6800
rect 67700 0 68100 6800
rect 84500 0 84900 6800
rect 101300 0 101700 6800
rect 118000 0 118500 6800
rect 119000 0 119600 6800
rect 211000 6892 211600 7300
rect 211000 0 211408 6892
rect 211500 0 212100 6800
rect 219700 0 220100 6800
rect 220700 0 221100 6800
rect 230700 0 231100 6800
rect 247500 0 247900 6800
rect 257500 0 257900 6800
rect 267500 0 267900 6800
rect 284300 0 284700 6800
rect 301100 0 301500 6800
rect 311100 0 311500 6800
rect 327900 0 328300 6800
rect 344700 0 345100 6800
rect 354700 0 355100 6800
rect 364700 0 365100 6800
rect 381500 0 381900 6800
rect 398300 0 398700 6800
rect 415100 0 415500 6800
rect 431900 0 432300 6800
rect 448700 0 449100 6800
rect 458700 0 459100 6800
rect 462700 0 463100 6800
rect 464700 0 465100 6800
rect 465900 0 466100 6800
rect 482700 0 483100 6800
<< psub >>
rect 97500 380826 97918 381244
rect 114300 380826 114718 381244
rect 131100 380826 131518 381244
rect 147900 380826 148318 381244
rect 204700 380826 205118 381244
rect 221500 380826 221918 381244
rect 248300 380826 248718 381244
rect 265100 380826 265518 381244
rect 281966 381134 282260 381164
rect 283544 381134 283838 381138
rect 281966 380948 282318 381134
rect 283494 380948 283838 381134
rect 281966 380826 282260 380948
rect 283544 380804 283838 380948
rect 47100 378426 47518 378844
rect 63900 378426 64318 378844
rect 91186 357820 315594 358080
rect 34450 145984 51252 146240
rect 120486 72030 120726 73098
<< subdiff >>
rect 91206 358040 315574 358060
rect 91206 357860 91226 358040
rect 315554 357860 315574 358040
rect 91206 357840 315574 357860
rect 120506 73058 120706 73078
rect 120506 72070 120526 73058
rect 120686 72070 120706 73058
rect 120506 72050 120706 72070
<< subdiffcont >>
rect 91226 357860 315554 358040
rect 120526 72070 120686 73058
<< mvsubdiff >>
rect 34470 146200 51232 146220
rect 34470 146024 34490 146200
rect 51212 146024 51232 146200
rect 34470 146004 51232 146024
<< mvsubdiffcont >>
rect 34490 146024 51212 146200
<< metal1 >>
rect 35168 392560 45584 405664
rect 51968 392560 62384 405664
rect 68768 392560 79184 405664
rect 85568 392560 95984 405664
rect 102368 392560 112784 405664
rect 119168 392560 129584 405664
rect 135968 392560 146384 405664
rect 192752 392560 203168 405664
rect 209552 392560 219968 405664
rect 236432 392560 246848 405664
rect 253232 392560 263648 405664
rect 269920 392560 280336 405664
rect 429296 392560 439824 405776
rect 446096 392560 456624 405776
rect 37520 381052 37632 381644
rect 33400 380580 34800 380600
rect 31939 380400 34800 380580
rect 31939 379588 33600 380400
rect 33400 379260 33600 379588
rect 31939 378268 33600 379260
rect 33400 377940 33600 378268
rect 31939 376948 33600 377940
rect 33400 376620 33600 376948
rect 31939 375628 33600 376620
rect 33400 375016 33600 375628
rect 31939 374024 33600 375016
rect 33400 373696 33600 374024
rect 31939 372704 33600 373696
rect 33400 372376 33600 372704
rect 31939 371384 33600 372376
rect 33400 370772 33600 371384
rect 31939 369780 33600 370772
rect 33400 369452 33600 369780
rect 31939 368460 33600 369452
rect 33400 368132 33600 368460
rect 31939 367140 33600 368132
rect 33400 366812 33600 367140
rect 31939 366000 33600 366812
rect 34600 366000 34800 380400
rect 37070 378686 37160 378696
rect 37070 378582 37160 378594
rect 37520 378686 37632 380996
rect 31939 365820 34800 366000
rect 33400 365800 34800 365820
rect 35550 378202 35872 378234
rect 35550 363800 35872 378058
rect 37050 378202 37182 378500
rect 37520 378494 37632 378594
rect 38192 381164 38304 381644
rect 38192 378660 38304 381108
rect 43008 380828 43120 381644
rect 44128 381388 44240 381644
rect 44128 381308 44240 381332
rect 43008 380732 43120 380772
rect 47712 380940 47824 381644
rect 47262 378686 47352 378702
rect 38192 378504 38304 378568
rect 38666 378660 38756 378670
rect 47262 378576 47352 378594
rect 47712 378686 47824 380884
rect 38666 378556 38756 378568
rect 47712 378544 47824 378594
rect 48384 381276 48496 381692
rect 48384 378660 48496 381220
rect 54320 380492 54432 381644
rect 53870 378686 53960 378696
rect 48384 378534 48496 378568
rect 48858 378660 48948 378676
rect 53870 378582 53960 378594
rect 54320 378686 54432 380436
rect 48858 378550 48948 378568
rect 54320 378536 54432 378594
rect 54992 380604 55104 381644
rect 54992 378660 55104 380548
rect 59808 380268 59920 381644
rect 60928 381388 61040 381644
rect 60928 381308 61040 381332
rect 59808 380188 59920 380212
rect 64512 380380 64624 381644
rect 64062 378686 64152 378702
rect 37050 378030 37182 378058
rect 38640 378202 38772 378478
rect 38640 378008 38772 378058
rect 47242 378202 47374 378515
rect 54992 378508 55104 378568
rect 55466 378660 55556 378670
rect 64062 378576 64152 378594
rect 64512 378686 64624 380324
rect 55466 378556 55556 378568
rect 64512 378556 64624 378594
rect 65184 380716 65296 381692
rect 65184 378660 65296 380660
rect 71120 379932 71232 381644
rect 70670 378686 70760 378696
rect 47242 378030 47374 378058
rect 48832 378202 48964 378493
rect 48832 378008 48964 378058
rect 53850 378202 53982 378500
rect 53850 378030 53982 378058
rect 55440 378202 55572 378478
rect 55440 378008 55572 378058
rect 64042 378202 64174 378515
rect 65184 378498 65296 378568
rect 65658 378660 65748 378676
rect 70670 378582 70760 378594
rect 71120 378686 71232 379876
rect 65658 378550 65748 378568
rect 71120 378540 71232 378594
rect 71792 380044 71904 381644
rect 71792 378660 71904 379988
rect 76608 379708 76720 381644
rect 77728 381388 77840 381644
rect 77728 381308 77840 381332
rect 76608 379612 76720 379652
rect 77110 380156 77228 380178
rect 76662 378686 76752 378702
rect 71792 378520 71904 378568
rect 72266 378660 72356 378670
rect 76662 378576 76752 378594
rect 77110 378686 77228 380100
rect 77110 378594 77112 378686
rect 77224 378594 77228 378686
rect 72266 378556 72356 378568
rect 77110 378554 77228 378594
rect 77784 379820 77898 379858
rect 77784 378660 77898 379764
rect 81312 379820 81424 381644
rect 81984 380156 82096 381692
rect 87470 381086 87560 381096
rect 87470 380982 87560 380994
rect 87920 381086 88032 381644
rect 87450 380602 87582 380900
rect 87450 380430 87582 380458
rect 81984 380060 82096 380100
rect 81312 379724 81424 379764
rect 87920 379372 88032 380994
rect 88592 381060 88704 381644
rect 88592 379484 88704 380968
rect 89066 381060 89156 381070
rect 89066 380956 89156 380968
rect 89040 380602 89172 380878
rect 89040 380408 89172 380458
rect 88592 379388 88704 379428
rect 87920 379276 88032 379316
rect 77896 378568 77898 378660
rect 77784 378534 77898 378568
rect 78258 378660 78348 378676
rect 78258 378550 78348 378568
rect 64042 378030 64174 378058
rect 65632 378202 65764 378493
rect 65632 378008 65764 378058
rect 70650 378202 70782 378500
rect 70650 378030 70782 378058
rect 72240 378202 72372 378478
rect 72240 378008 72372 378058
rect 76642 378202 76774 378515
rect 76642 378030 76774 378058
rect 78232 378202 78364 378493
rect 78232 378008 78364 378058
rect 93380 374927 93436 381644
rect 94528 381388 94640 381644
rect 94528 381308 94640 381332
rect 97662 381086 97752 381102
rect 97662 380976 97752 380994
rect 98112 381086 98224 381644
rect 97642 380602 97774 380915
rect 97642 380430 97774 380458
rect 98112 379260 98224 380994
rect 98784 381060 98896 381692
rect 104270 381086 104360 381096
rect 98784 379596 98896 380968
rect 99258 381060 99348 381076
rect 104270 380982 104360 380994
rect 104720 381086 104832 381644
rect 99258 380950 99348 380968
rect 99232 380602 99364 380893
rect 99232 380408 99364 380458
rect 104250 380602 104382 380900
rect 104250 380430 104382 380458
rect 98784 379500 98896 379540
rect 98112 379164 98224 379204
rect 104720 378924 104832 380994
rect 105392 381060 105504 381644
rect 105392 379036 105504 380968
rect 105866 381060 105956 381070
rect 105866 380956 105956 380968
rect 105840 380602 105972 380878
rect 105840 380408 105972 380458
rect 105392 378961 105504 378980
rect 104720 378843 104832 378868
rect 93380 374192 93436 374257
rect 110180 374927 110236 381692
rect 111328 381388 111440 381644
rect 111328 381308 111440 381332
rect 114462 381086 114552 381102
rect 114462 380976 114552 380994
rect 114912 381086 115024 381644
rect 114442 380602 114574 380915
rect 114442 380430 114574 380458
rect 114912 378812 115024 380994
rect 115584 381060 115696 381692
rect 121070 381086 121160 381096
rect 115584 379148 115696 380968
rect 116058 381060 116148 381076
rect 121070 380982 121160 380994
rect 121520 381086 121632 381644
rect 116058 380950 116148 380968
rect 116032 380602 116164 380893
rect 116032 380408 116164 380458
rect 121050 380602 121182 380900
rect 121050 380430 121182 380458
rect 115584 379052 115696 379092
rect 114912 378716 115024 378756
rect 121520 378476 121632 380994
rect 122192 381060 122304 381644
rect 122192 378588 122304 380968
rect 122666 381060 122756 381070
rect 122666 380956 122756 380968
rect 122640 380602 122772 380878
rect 122640 380408 122772 380458
rect 122192 378492 122304 378532
rect 121520 378380 121632 378420
rect 110180 374192 110236 374257
rect 126980 374927 127036 381692
rect 128128 381388 128240 381644
rect 128128 381308 128240 381332
rect 131262 381086 131352 381102
rect 131262 380976 131352 380994
rect 131712 381086 131824 381644
rect 131242 380602 131374 380915
rect 131242 380430 131374 380458
rect 131712 378364 131824 380994
rect 132384 381060 132496 381692
rect 137870 381086 137960 381096
rect 132384 378700 132496 380968
rect 132858 381060 132948 381076
rect 137870 380982 137960 380994
rect 138320 381086 138432 381644
rect 132858 380950 132948 380968
rect 132832 380602 132964 380893
rect 132832 380408 132964 380458
rect 137850 380602 137982 380900
rect 137850 380430 137982 380458
rect 132384 378604 132496 378644
rect 131712 378268 131824 378308
rect 138320 378028 138432 380994
rect 138992 381060 139104 381644
rect 138992 378140 139104 380968
rect 139466 381060 139556 381070
rect 139466 380956 139556 380968
rect 139440 380602 139572 380878
rect 139440 380408 139572 380458
rect 138992 378044 139104 378084
rect 138320 377932 138432 377972
rect 126980 374192 127036 374257
rect 143780 374927 143836 381692
rect 144928 381388 145040 381644
rect 144928 381308 145040 381332
rect 148062 381086 148152 381102
rect 148062 380976 148152 380994
rect 148512 381086 148624 381644
rect 148042 380602 148174 380915
rect 148042 380430 148174 380458
rect 148512 377916 148624 380994
rect 149184 381060 149296 381692
rect 194670 381086 194760 381096
rect 149184 378252 149296 380968
rect 149658 381060 149748 381076
rect 194670 380982 194760 380994
rect 195120 381086 195232 381644
rect 149658 380950 149748 380968
rect 149632 380602 149764 380893
rect 149632 380408 149764 380458
rect 194650 380602 194782 380900
rect 194650 380430 194782 380458
rect 149184 378156 149296 378196
rect 148512 377820 148624 377860
rect 195120 377580 195232 380994
rect 195792 381060 195904 381644
rect 195792 377692 195904 380968
rect 196266 381060 196356 381070
rect 196266 380956 196356 380968
rect 196240 380602 196372 380878
rect 196240 380408 196372 380458
rect 195792 377596 195904 377636
rect 195120 377484 195232 377524
rect 143780 374192 143836 374257
rect 200580 374927 200636 381692
rect 201712 381388 201824 381644
rect 201712 381308 201824 381332
rect 204862 381086 204952 381102
rect 204862 380976 204952 380994
rect 205312 381086 205424 381644
rect 204842 380602 204974 380915
rect 204842 380430 204974 380458
rect 205312 377468 205424 380994
rect 205984 381060 206096 381692
rect 211470 381086 211560 381096
rect 205984 377804 206096 380968
rect 206458 381060 206548 381076
rect 211470 380982 211560 380994
rect 211920 381086 212032 381644
rect 206458 380950 206548 380968
rect 206432 380602 206564 380893
rect 206432 380408 206564 380458
rect 211450 380602 211582 380900
rect 211450 380430 211582 380458
rect 205984 377708 206096 377748
rect 205312 377372 205424 377412
rect 211920 377132 212032 380994
rect 212592 381060 212704 381644
rect 212592 377244 212704 380968
rect 213066 381060 213156 381070
rect 213066 380956 213156 380968
rect 213040 380602 213172 380878
rect 213040 380408 213172 380458
rect 212592 377148 212704 377188
rect 211920 377036 212032 377076
rect 200580 374192 200636 374257
rect 217380 374927 217436 381692
rect 218512 381388 218624 381644
rect 218512 381308 218624 381332
rect 221662 381086 221752 381102
rect 221662 380976 221752 380994
rect 222112 381086 222224 381644
rect 221642 380602 221774 380915
rect 221642 380430 221774 380458
rect 222112 377020 222224 380994
rect 222784 381060 222896 381692
rect 238270 381086 238360 381096
rect 222784 377356 222896 380968
rect 223258 381060 223348 381076
rect 238270 380982 238360 380994
rect 238720 381086 238832 381644
rect 223258 380950 223348 380968
rect 223232 380602 223364 380893
rect 223232 380408 223364 380458
rect 238250 380602 238382 380900
rect 238250 380430 238382 380458
rect 222784 377260 222896 377300
rect 222112 376924 222224 376964
rect 238720 376684 238832 380994
rect 239392 381060 239504 381644
rect 239392 376796 239504 380968
rect 239866 381060 239956 381070
rect 239866 380956 239956 380968
rect 239840 380602 239972 380878
rect 239840 380408 239972 380458
rect 239392 376700 239504 376740
rect 238720 376588 238832 376628
rect 217380 374192 217436 374257
rect 244180 374927 244236 381692
rect 245280 381388 245392 381644
rect 245280 381308 245392 381332
rect 248462 381086 248552 381102
rect 248462 380976 248552 380994
rect 248912 381086 249024 381644
rect 248442 380602 248574 380915
rect 248442 380430 248574 380458
rect 248912 376572 249024 380994
rect 249584 381060 249696 381692
rect 255070 381086 255160 381096
rect 249584 376908 249696 380968
rect 250058 381060 250148 381076
rect 255070 380982 255160 380994
rect 255520 381086 255632 381644
rect 250058 380950 250148 380968
rect 250032 380602 250164 380893
rect 250032 380408 250164 380458
rect 255050 380602 255182 380900
rect 255050 380430 255182 380458
rect 249584 376812 249696 376852
rect 248912 376476 249024 376516
rect 255520 376236 255632 380994
rect 256192 381060 256304 381644
rect 256192 376348 256304 380968
rect 256666 381060 256756 381070
rect 256666 380956 256756 380968
rect 256640 380602 256772 380878
rect 256640 380408 256772 380458
rect 256192 376252 256304 376292
rect 255520 376140 255632 376180
rect 244180 374192 244236 374257
rect 260980 374927 261036 381692
rect 262080 381388 262192 381644
rect 262080 381308 262192 381332
rect 265262 381086 265352 381102
rect 265262 380976 265352 380994
rect 265712 381086 265824 381644
rect 265242 380602 265374 380915
rect 265242 380430 265374 380458
rect 265712 376124 265824 380994
rect 266384 381060 266496 381692
rect 271870 381086 271960 381096
rect 266384 376460 266496 380968
rect 266858 381060 266948 381076
rect 271870 380982 271960 380994
rect 272320 381086 272432 381644
rect 266858 380950 266948 380968
rect 266832 380602 266964 380893
rect 266832 380408 266964 380458
rect 271850 380602 271982 380900
rect 271850 380430 271982 380458
rect 266384 376364 266496 376404
rect 265712 376028 265824 376068
rect 272320 375788 272432 380994
rect 272992 381060 273104 381644
rect 272992 375900 273104 380968
rect 273466 381060 273556 381070
rect 273466 380956 273556 380968
rect 273440 380602 273572 380878
rect 273440 380408 273572 380458
rect 272992 375804 273104 375844
rect 272320 375692 272432 375732
rect 260980 374192 261036 374257
rect 277780 374927 277836 381692
rect 278880 381388 278992 381644
rect 278880 381308 278992 381332
rect 281966 381155 282260 381164
rect 281966 380915 281989 381155
rect 282229 381134 282260 381155
rect 282062 381086 282152 381102
rect 282062 380976 282152 380994
rect 282229 380948 282275 381134
rect 282512 381086 282624 381644
rect 282229 380915 282260 380948
rect 281966 380869 282260 380915
rect 282042 380602 282174 380869
rect 282042 380430 282174 380458
rect 282512 375676 282624 380994
rect 283184 381060 283296 381692
rect 283544 381134 283838 381138
rect 283184 376012 283296 380968
rect 283537 381133 283838 381134
rect 283537 380948 283583 381133
rect 283658 381060 283748 381076
rect 283658 380950 283748 380968
rect 283544 380893 283583 380948
rect 283823 380893 283838 381133
rect 283544 380847 283838 380893
rect 283632 380602 283764 380847
rect 283632 380408 283764 380458
rect 427220 376000 428212 381616
rect 428540 376000 429532 381616
rect 429860 376000 430852 381616
rect 431180 376000 432172 381616
rect 432784 376000 433776 381616
rect 434104 376000 435096 381616
rect 435424 376000 436416 381616
rect 437028 376000 438020 381616
rect 438348 376000 439340 381616
rect 439668 376000 440660 381616
rect 440988 376000 441980 381616
rect 444020 376000 445012 381659
rect 445340 376000 446332 381659
rect 446660 376000 447652 381659
rect 447980 376000 448972 381659
rect 449584 376000 450576 381659
rect 450904 376000 451896 381659
rect 452224 376000 453216 381659
rect 453828 376000 454820 381659
rect 455148 376000 456140 381659
rect 456468 376000 457460 381659
rect 457788 376000 458780 381659
rect 466820 376000 467812 381639
rect 468140 376000 469132 381639
rect 469460 376000 470452 381639
rect 470780 376000 471772 381639
rect 472384 376000 473376 381639
rect 473704 376000 474696 381639
rect 475024 376000 476016 381639
rect 476628 376000 477620 381639
rect 477948 376000 478940 381639
rect 479268 376000 480260 381639
rect 480588 376000 481580 381639
rect 283184 375916 283296 375956
rect 282512 375580 282624 375620
rect 427200 375800 442000 376000
rect 277780 374192 277836 374257
rect 427200 374200 427400 375800
rect 441800 374200 442000 375800
rect 427200 374000 442000 374200
rect 444000 375800 458800 376000
rect 444000 374200 444200 375800
rect 458600 374200 458800 375800
rect 444000 374000 458800 374200
rect 466800 375800 481600 376000
rect 466800 374200 467000 375800
rect 481400 374200 481600 375800
rect 466800 374000 481600 374200
rect 466820 373968 467812 374000
rect 468140 373968 469132 374000
rect 469460 373968 470452 374000
rect 470780 373968 471772 374000
rect 472384 373968 473376 374000
rect 473704 373968 474696 374000
rect 475024 373968 476016 374000
rect 476628 373968 477620 374000
rect 477948 373968 478940 374000
rect 479268 373968 480260 374000
rect 480588 373968 481580 374000
rect 471400 373500 472100 373600
rect 471400 373400 471500 373500
rect 470759 373000 471500 373400
rect 472000 373000 472100 373500
rect 471400 372900 472100 373000
rect 480624 370514 480662 370636
rect 480718 370514 482640 370636
rect 481824 369264 481908 369376
rect 481964 369264 482608 369376
rect 493584 367920 506688 378448
rect 33400 363780 35872 363800
rect 31949 363600 35872 363780
rect 31949 362788 33600 363600
rect 33400 362460 33600 362788
rect 31949 361468 33600 362460
rect 33400 361140 33600 361468
rect 31949 360148 33600 361140
rect 33400 359820 33600 360148
rect 31949 358828 33600 359820
rect 33400 358216 33600 358828
rect 31949 357224 33600 358216
rect 33400 356896 33600 357224
rect 31949 355904 33600 356896
rect 33400 355576 33600 355904
rect 31949 354584 33600 355576
rect 33400 353972 33600 354584
rect 31949 352980 33600 353972
rect 33400 352652 33600 352980
rect 31949 351660 33600 352652
rect 33400 351332 33600 351660
rect 31949 350340 33600 351332
rect 33400 350012 33600 350340
rect 31949 349200 33600 350012
rect 34600 363201 35872 363600
rect 63378 367542 64890 367668
rect 63378 366912 63504 367542
rect 64764 366912 64890 367542
rect 63378 366786 64890 366912
rect 34600 349200 34800 363201
rect 63378 360486 63756 366786
rect 320670 365486 322812 365612
rect 320670 364604 320796 365486
rect 322686 364604 322812 365486
rect 320670 364478 322812 364604
rect 320670 363512 321048 364478
rect 328700 364100 329100 364880
rect 328500 364000 329300 364100
rect 319127 363388 321057 363512
rect 328500 363400 328600 364000
rect 329200 363400 329300 364000
rect 66024 361620 66906 361746
rect 65268 360864 65772 360990
rect 65268 360418 65394 360864
rect 65016 360360 65394 360418
rect 65646 360360 65772 360864
rect 65016 360294 65772 360360
rect 65268 360234 65772 360294
rect 66024 360360 66150 361620
rect 66780 360360 66906 361620
rect 319127 361130 319251 363388
rect 320670 363384 321048 363388
rect 328500 363300 329300 363400
rect 472400 363780 478000 363800
rect 472400 363600 482652 363780
rect 321048 362502 323442 362628
rect 321048 361998 322056 362502
rect 321048 361746 321426 361998
rect 321930 361872 322056 361998
rect 323316 361872 323442 362502
rect 321930 361746 323442 361872
rect 334336 362400 339936 362949
rect 340548 362400 346148 362949
rect 334336 362200 346200 362400
rect 316764 360990 317772 361116
rect 319127 361006 319548 361130
rect 316764 360612 316890 360990
rect 317646 360960 317772 360990
rect 317646 360800 319742 360960
rect 334336 360800 334600 362200
rect 346000 360800 346200 362200
rect 317646 360612 317772 360800
rect 316764 360486 317772 360612
rect 334336 360600 346200 360800
rect 66024 360234 66906 360360
rect 64762 360116 64778 360172
rect 64940 360116 64956 360172
rect 66070 359728 66230 360234
rect 64936 359568 66230 359728
rect 63000 358880 63630 359040
rect 63000 358470 63504 358880
rect 63000 358092 63126 358470
rect 63378 358092 63504 358470
rect 63644 358418 63662 358494
rect 63798 358418 63812 358494
rect 64316 358418 64332 358494
rect 64472 358418 64484 358494
rect 66070 358144 66230 359568
rect 63000 357966 63504 358092
rect 64800 357984 66230 358144
rect 148820 356852 149276 357860
rect 272636 357648 272692 357664
rect 272636 357360 272692 357390
rect 272888 357648 272944 357664
rect 272888 357360 272944 357390
rect 273140 357648 273196 357664
rect 273140 357360 273196 357390
rect 273392 357648 273448 357664
rect 273392 357360 273448 357390
rect 273644 357648 273700 357664
rect 273644 357360 273700 357390
rect 273896 357648 273952 357664
rect 273896 357360 273952 357390
rect 274148 357648 274204 357664
rect 274148 357360 274204 357390
rect 89798 356090 89824 356146
rect 90170 356090 90192 356146
rect 89798 355846 89824 355902
rect 90170 355846 90192 355902
rect 89798 355602 89824 355658
rect 90170 355602 90192 355658
rect 89798 355358 89824 355414
rect 90170 355358 90192 355414
rect 89798 355114 89824 355170
rect 90170 355114 90192 355170
rect 89798 354870 89824 354926
rect 90170 354870 90192 354926
rect 89798 354626 89824 354682
rect 90170 354626 90192 354682
rect 89798 354382 89824 354438
rect 90170 354382 90192 354438
rect 89798 354138 89824 354194
rect 90170 354138 90192 354194
rect 89798 353894 89824 353950
rect 90170 353894 90192 353950
rect 31949 349020 34800 349200
rect 33400 349000 34800 349020
rect 472400 349200 472600 363600
rect 477800 362788 482652 363600
rect 477800 362460 478000 362788
rect 477800 361468 482652 362460
rect 477800 361140 478000 361468
rect 477800 360148 482652 361140
rect 477800 359820 478000 360148
rect 477800 358828 482652 359820
rect 477800 358216 478000 358828
rect 477800 357224 482652 358216
rect 477800 356896 478000 357224
rect 477800 355904 482652 356896
rect 477800 355576 478000 355904
rect 477800 354584 482652 355576
rect 477800 353972 478000 354584
rect 477800 352980 482652 353972
rect 477800 352652 478000 352980
rect 477800 351660 482652 352652
rect 477800 351332 478000 351660
rect 477800 350340 482652 351332
rect 493584 351120 506688 361648
rect 477800 350012 478000 350340
rect 477800 349200 482652 350012
rect 472400 349020 482652 349200
rect 472400 349000 478000 349020
rect 410130 341712 412020 342972
rect 410130 340578 410256 341712
rect 411894 340578 412020 341712
rect 410130 340452 412020 340578
rect 32792 338042 32808 338132
rect 32900 338042 32918 338132
rect 32975 338016 33226 338148
rect 33370 338016 33420 338148
rect 31908 337568 32808 337680
rect 32900 337568 34020 337680
rect 34076 337568 34116 337680
rect 31908 337008 32782 337120
rect 32874 337008 34356 337120
rect 34412 337008 34452 337120
rect 32766 336558 32782 336648
rect 32874 336558 32892 336648
rect 32953 336538 33226 336670
rect 33370 336538 33398 336670
rect 7840 324352 20944 334880
rect 493584 334320 506688 344848
rect 31920 333312 32228 333424
rect 32284 333312 32368 333424
rect 477520 332418 477548 332524
rect 477644 332418 477656 332524
rect 477712 332400 477862 332528
rect 477984 332400 478004 332528
rect 31908 332192 34468 332304
rect 34524 332192 34564 332304
rect 477502 332080 477548 332192
rect 477644 332080 482160 332192
rect 482216 332080 482608 332192
rect 477531 331474 477552 331596
rect 477648 331474 481166 331596
rect 481222 331474 482640 331596
rect 477538 330986 477552 331092
rect 477648 330986 477674 331092
rect 477736 330976 477862 331104
rect 477984 330976 478006 331104
rect 32792 327850 32808 327940
rect 32900 327850 32918 327940
rect 32975 327824 33226 327956
rect 33370 327824 33414 327956
rect 31908 327376 32808 327488
rect 32900 327376 34132 327488
rect 34188 327376 34228 327488
rect 31908 326704 32782 326816
rect 32874 326704 34244 326816
rect 34300 326704 34340 326816
rect 32766 326254 32782 326344
rect 32874 326254 32892 326344
rect 32953 326234 33226 326366
rect 33370 326234 33398 326366
rect 32792 321242 32808 321332
rect 32900 321242 32918 321332
rect 32975 321216 33226 321348
rect 33370 321216 33414 321348
rect 31908 320768 32808 320880
rect 32900 320768 33460 320880
rect 33516 320768 33576 320880
rect 31908 320208 32782 320320
rect 32874 320208 33796 320320
rect 33852 320208 33892 320320
rect 32766 319758 32782 319848
rect 32874 319758 32892 319848
rect 32953 319738 33226 319870
rect 33370 319738 33398 319870
rect 7840 307552 20944 318080
rect 493584 317520 506688 328048
rect 332990 316862 333046 316887
rect 31920 316512 32228 316624
rect 32284 316512 32368 316624
rect 332990 316440 333046 316684
rect 333368 316862 333424 316887
rect 333368 316440 333424 316684
rect 333872 316862 333928 316887
rect 333872 316440 333928 316684
rect 336644 316862 336700 316887
rect 336644 316440 336700 316684
rect 337148 316862 337204 316887
rect 337148 316440 337204 316684
rect 337652 316862 337708 316887
rect 337652 316440 337708 316684
rect 340424 316862 340480 316887
rect 340424 316440 340480 316684
rect 340928 316862 340984 316887
rect 340928 316440 340984 316684
rect 341432 316862 341488 316887
rect 341432 316440 341488 316684
rect 344204 316862 344260 316887
rect 344204 316440 344260 316684
rect 344708 316862 344764 316887
rect 344708 316440 344764 316684
rect 345212 316862 345268 316887
rect 345212 316440 345268 316684
rect 347984 316862 348040 316887
rect 347984 316440 348040 316684
rect 348488 316862 348544 316887
rect 348488 316440 348544 316684
rect 348992 316862 349048 316887
rect 348992 316440 349048 316684
rect 351764 316862 351820 316887
rect 351764 316440 351820 316684
rect 352268 316862 352324 316887
rect 352268 316440 352324 316684
rect 352772 316862 352828 316887
rect 352772 316440 352828 316684
rect 355544 316862 355600 316887
rect 355544 316440 355600 316684
rect 356048 316862 356104 316887
rect 356048 316440 356104 316684
rect 356552 316862 356608 316887
rect 356552 316440 356608 316684
rect 359324 316862 359380 316887
rect 359324 316440 359380 316684
rect 359828 316862 359884 316887
rect 359828 316440 359884 316684
rect 360332 316862 360388 316887
rect 360332 316440 360388 316684
rect 363104 316862 363160 316887
rect 363104 316440 363160 316684
rect 363608 316862 363664 316887
rect 363608 316440 363664 316684
rect 364112 316862 364168 316887
rect 364112 316440 364168 316684
rect 366758 316862 366814 316887
rect 366758 316440 366814 316684
rect 367262 316862 367318 316887
rect 367262 316440 367318 316684
rect 367766 316862 367822 316887
rect 367766 316440 367822 316684
rect 370538 316862 370594 316887
rect 370538 316440 370594 316684
rect 371042 316862 371098 316887
rect 371042 316440 371098 316684
rect 371546 316862 371602 316887
rect 371546 316440 371602 316684
rect 374318 316862 374374 316887
rect 374318 316440 374374 316684
rect 374822 316862 374878 316887
rect 374822 316440 374878 316684
rect 375326 316862 375382 316887
rect 375326 316440 375382 316684
rect 378098 316862 378154 316887
rect 378098 316440 378154 316684
rect 378602 316862 378658 316887
rect 378602 316440 378658 316684
rect 379106 316862 379162 316887
rect 379106 316440 379162 316684
rect 381878 316862 381934 316887
rect 381878 316440 381934 316684
rect 382382 316862 382438 316887
rect 382382 316440 382438 316684
rect 382886 316862 382942 316887
rect 382886 316440 382942 316684
rect 385658 316862 385714 316887
rect 385658 316440 385714 316684
rect 386162 316862 386218 316887
rect 386162 316440 386218 316684
rect 386666 316862 386722 316887
rect 386666 316440 386722 316684
rect 389438 316862 389494 316887
rect 389438 316440 389494 316684
rect 389942 316862 389998 316887
rect 389942 316440 389998 316684
rect 390446 316862 390502 316887
rect 390446 316440 390502 316684
rect 395612 316862 395668 316887
rect 395612 316440 395668 316684
rect 396116 316862 396172 316887
rect 396116 316440 396172 316684
rect 396872 316862 396928 316887
rect 396872 316440 396928 316684
rect 398006 316862 398062 316887
rect 398006 316496 398062 316684
rect 401534 316862 401590 316887
rect 401534 316440 401590 316684
rect 402038 316862 402094 316887
rect 402038 316440 402094 316684
rect 402542 316862 402598 316887
rect 402542 316440 402598 316684
rect 403046 316862 403102 316887
rect 403046 316440 403102 316684
rect 403550 316862 403606 316887
rect 403550 316440 403606 316684
rect 404054 316862 404110 316887
rect 404054 316440 404110 316684
rect 404558 316862 404614 316887
rect 404558 316440 404614 316684
rect 405062 316862 405118 316887
rect 405062 316440 405118 316684
rect 405566 316862 405622 316887
rect 405566 316440 405622 316684
rect 406070 316862 406126 316887
rect 406070 316440 406126 316684
rect 408842 316862 408898 316887
rect 408842 316440 408898 316684
rect 409346 316862 409402 316887
rect 409346 316440 409402 316684
rect 409850 316862 409906 316887
rect 409850 316440 409906 316684
rect 412622 316862 412678 316887
rect 412622 316440 412678 316684
rect 413126 316862 413182 316887
rect 413126 316440 413182 316684
rect 413630 316862 413686 316887
rect 413630 316440 413686 316684
rect 416402 316862 416458 316887
rect 416402 316440 416458 316684
rect 416906 316862 416962 316887
rect 416906 316440 416962 316684
rect 417410 316862 417466 316887
rect 417410 316440 417466 316684
rect 420182 316862 420238 316887
rect 420182 316440 420238 316684
rect 420686 316862 420742 316887
rect 420686 316440 420742 316684
rect 421190 316862 421246 316887
rect 421190 316440 421246 316684
rect 423962 316862 424018 316887
rect 423962 316440 424018 316684
rect 424466 316862 424522 316887
rect 424466 316440 424522 316684
rect 424970 316862 425026 316887
rect 424970 316440 425026 316684
rect 427616 316862 427672 316887
rect 427616 316440 427672 316684
rect 428120 316862 428176 316887
rect 428120 316440 428176 316684
rect 428624 316862 428680 316887
rect 428624 316440 428680 316684
rect 431396 316862 431452 316887
rect 431396 316440 431452 316684
rect 431900 316862 431956 316887
rect 431900 316440 431956 316684
rect 432404 316862 432460 316887
rect 432404 316440 432460 316684
rect 435176 316862 435232 316887
rect 435176 316440 435232 316684
rect 435680 316862 435736 316887
rect 435680 316440 435736 316684
rect 436184 316862 436240 316887
rect 436184 316440 436240 316684
rect 438956 316862 439012 316887
rect 438956 316440 439012 316684
rect 439460 316862 439516 316887
rect 439460 316440 439516 316684
rect 439964 316862 440020 316887
rect 439964 316440 440020 316684
rect 442736 316862 442792 316887
rect 442736 316440 442792 316684
rect 443240 316862 443296 316887
rect 443240 316440 443296 316684
rect 443744 316862 443800 316887
rect 443744 316440 443800 316684
rect 446516 316862 446572 316887
rect 446516 316440 446572 316684
rect 447020 316862 447076 316887
rect 447020 316440 447076 316684
rect 447524 316862 447580 316887
rect 447524 316440 447580 316684
rect 450296 316862 450352 316887
rect 450296 316440 450352 316684
rect 450800 316862 450856 316887
rect 450800 316440 450856 316684
rect 451304 316862 451360 316887
rect 451304 316440 451360 316684
rect 454076 316862 454132 316887
rect 454076 316440 454132 316684
rect 454580 316862 454636 316887
rect 454580 316440 454636 316684
rect 455084 316862 455140 316887
rect 455084 316440 455140 316684
rect 457730 316862 457786 316887
rect 457730 316440 457786 316684
rect 458234 316862 458290 316887
rect 458234 316440 458290 316684
rect 458738 316862 458794 316887
rect 458738 316440 458794 316684
rect 461510 316862 461566 316887
rect 461510 316440 461566 316684
rect 462014 316862 462070 316887
rect 462014 316440 462070 316684
rect 462518 316862 462574 316887
rect 462518 316440 462574 316684
rect 465290 316862 465346 316887
rect 465290 316440 465346 316684
rect 465794 316862 465850 316887
rect 465794 316440 465850 316684
rect 466298 316862 466354 316887
rect 466298 316440 466354 316684
rect 477520 315618 477548 315724
rect 477644 315618 477656 315724
rect 477712 315600 477862 315728
rect 477984 315600 478004 315728
rect 31908 315392 33908 315504
rect 33964 315392 34004 315504
rect 477502 315280 477548 315392
rect 477644 315280 482160 315392
rect 482216 315280 482608 315392
rect 477997 314796 481418 314882
rect 477531 314674 477552 314796
rect 477648 314760 481418 314796
rect 481474 314760 482640 314882
rect 477648 314674 478114 314760
rect 477538 314186 477552 314292
rect 477648 314186 477674 314292
rect 477736 314176 477862 314304
rect 477984 314176 478006 314304
rect 42714 314092 43344 314118
rect 40606 313892 47857 314092
rect 35028 313488 36540 313614
rect 35028 312984 35154 313488
rect 35910 313362 36540 313488
rect 38396 313604 38596 313616
rect 35910 312984 36036 313362
rect 38396 313329 38413 313604
rect 38578 313329 38596 313604
rect 38396 313314 38596 313329
rect 39872 313597 40072 313616
rect 39872 313333 39889 313597
rect 40051 313333 40072 313597
rect 40606 313388 40806 313892
rect 41725 313623 41985 313646
rect 41725 313438 41744 313623
rect 41962 313438 41985 313623
rect 41725 313338 41985 313438
rect 42714 313614 43344 313892
rect 39872 313314 40072 313333
rect 35028 312858 36036 312984
rect 42714 312858 42840 313614
rect 43218 312858 43344 313614
rect 45447 313601 45647 313624
rect 45447 313339 45467 313601
rect 45631 313339 45647 313601
rect 45447 313322 45647 313339
rect 46923 313610 47123 313624
rect 46923 313336 46935 313610
rect 47111 313336 47123 313610
rect 47657 313388 47857 313892
rect 48764 313634 49026 313649
rect 48764 313456 48779 313634
rect 49011 313456 49026 313634
rect 48764 313345 49026 313456
rect 60228 313456 61362 313488
rect 60228 313362 62712 313456
rect 46923 313322 47123 313336
rect 60228 313110 60354 313362
rect 61236 313296 62712 313362
rect 61236 313110 61362 313296
rect 60228 312984 61362 313110
rect 42714 312732 43344 312858
rect 64386 312732 65520 312858
rect 64386 312580 64512 312732
rect 59498 312480 64512 312580
rect 65394 312480 65520 312732
rect 59498 312380 65520 312480
rect 59498 312160 59698 312380
rect 64386 312354 65520 312380
rect 56900 311960 59698 312160
rect 60228 311891 61362 311976
rect 60228 311850 62828 311891
rect 48888 311442 51408 311472
rect 32792 311050 32808 311140
rect 32900 311050 32918 311140
rect 32975 311024 33226 311156
rect 33370 311024 33414 311156
rect 41674 311122 43626 311434
rect 48725 311130 51408 311442
rect 60228 311278 60354 311850
rect 42714 310842 43344 310968
rect 31908 310576 32808 310688
rect 32900 310576 33572 310688
rect 33628 310576 33668 310688
rect 42714 310338 42840 310842
rect 43218 310338 43344 310842
rect 42714 310212 43344 310338
rect 49896 310842 50526 310968
rect 49896 310338 50022 310842
rect 50400 310338 50526 310842
rect 49896 310212 50526 310338
rect 31908 309904 32782 310016
rect 32874 309904 33684 310016
rect 33740 309904 33780 310016
rect 32766 309454 32782 309544
rect 32874 309454 32892 309544
rect 32953 309434 33226 309566
rect 33370 309434 33398 309566
rect 42866 309544 43066 310212
rect 50048 309552 50248 310212
rect 50904 309708 51408 311130
rect 56896 311220 60354 311278
rect 61236 311731 62828 311850
rect 61236 311220 61362 311731
rect 56896 311078 61362 311220
rect 68544 311220 69552 311346
rect 68544 310995 68670 311220
rect 67708 310968 68670 310995
rect 69426 310968 69552 311220
rect 67708 310842 69552 310968
rect 67708 310835 69380 310842
rect 52672 310398 52708 310598
rect 52947 310398 54094 310598
rect 57886 310424 58126 310447
rect 57886 310414 57903 310424
rect 41732 309344 43066 309544
rect 48849 309352 50248 309552
rect 50526 309582 51408 309708
rect 50526 309078 50652 309582
rect 51282 309078 51408 309582
rect 50526 308952 51408 309078
rect 53900 308560 54100 310300
rect 56898 310214 57903 310414
rect 57886 310206 57903 310214
rect 58105 310414 58126 310424
rect 58105 310214 68976 310414
rect 69088 310214 69188 310414
rect 58105 310206 58126 310214
rect 57886 310183 58126 310206
rect 58464 309582 58968 309708
rect 58464 309468 58590 309582
rect 56904 309268 58590 309468
rect 58464 308952 58590 309268
rect 58842 308952 58968 309582
rect 58464 308826 58968 308952
rect 53900 308439 54100 308460
rect 32344 304430 32358 304556
rect 32430 304430 32442 304556
rect 32528 304462 32566 304526
rect 32632 304462 32666 304526
rect 31908 303968 32566 304080
rect 32632 303968 32900 304080
rect 32956 303968 32996 304080
rect 31908 303408 32540 303520
rect 32612 303408 33236 303520
rect 33292 303408 33332 303520
rect 32340 302836 32358 302962
rect 32512 302860 32540 302936
rect 32612 302860 32644 302936
rect 7840 290752 20944 301280
rect 493584 300720 506688 311248
rect 31920 299712 32228 299824
rect 32284 299712 32368 299824
rect 477520 298818 477548 298924
rect 477644 298818 477656 298924
rect 477712 298800 477862 298928
rect 477984 298800 478004 298928
rect 31908 298592 33348 298704
rect 33404 298592 33444 298704
rect 477965 298592 481670 298656
rect 477502 298480 477548 298592
rect 477644 298534 481670 298592
rect 481726 298534 482640 298656
rect 477644 298480 478114 298534
rect 477955 297996 480914 298046
rect 477531 297874 477552 297996
rect 477648 297924 480914 297996
rect 480970 297924 482640 298046
rect 477648 297874 478114 297924
rect 477538 297386 477552 297492
rect 477648 297386 477674 297492
rect 477736 297376 477862 297504
rect 477984 297376 478006 297504
rect 32346 294118 32358 294244
rect 32532 294140 32562 294224
rect 32630 294140 32662 294224
rect 31908 293776 32562 293888
rect 32630 293776 33012 293888
rect 33068 293776 33108 293888
rect 31908 293104 32540 293216
rect 32610 293104 33124 293216
rect 33180 293104 33220 293216
rect 32332 292524 32358 292650
rect 32508 292546 32540 292630
rect 32610 292546 32638 292630
rect 32330 288570 32358 288694
rect 32454 288570 32490 288694
rect 32546 288596 32570 288670
rect 32656 288596 32678 288670
rect 32094 288270 32108 288326
rect 32164 288270 32570 288326
rect 32656 288270 32674 288326
rect 32344 287776 32358 287904
rect 32528 287804 32554 287882
rect 32628 287804 32660 287882
rect 31920 287168 32108 287280
rect 32164 287168 32340 287280
rect 32396 287168 32436 287280
rect 31920 286608 32554 286720
rect 32628 286608 32676 286720
rect 32732 286608 32772 286720
rect 7840 273840 20944 284368
rect 31920 282912 32228 283024
rect 32284 282912 32368 283024
rect 31920 281792 32788 281904
rect 32844 281792 32884 281904
rect 33092 277450 33108 277540
rect 33200 277450 33218 277540
rect 33275 277424 33526 277556
rect 33670 277424 33714 277556
rect 31920 276976 32452 277088
rect 32508 276976 33108 277088
rect 33200 276976 33234 277088
rect 31920 276304 32564 276416
rect 32620 276304 33082 276416
rect 33174 276304 33210 276416
rect 33066 275854 33082 275944
rect 33174 275854 33192 275944
rect 33253 275834 33526 275966
rect 33670 275834 33698 275966
rect 33695 257206 34047 257276
rect 33695 257144 33739 257206
rect 31908 256496 33739 257144
rect 33695 255980 33739 256496
rect 31908 255332 33739 255980
rect 7840 244720 20944 255248
rect 33695 254701 33739 255332
rect 31908 254062 33739 254701
rect 33994 254062 34047 257206
rect 31908 254053 34047 254062
rect 33695 254010 34047 254053
rect 478860 246440 478898 246562
rect 478954 246440 482640 246562
rect 481824 245280 481908 245392
rect 481964 245280 482608 245392
rect 63756 244692 64764 244818
rect 63756 243936 63882 244692
rect 64638 243936 64764 244692
rect 493584 243936 506688 254464
rect 63756 243882 64764 243936
rect 67158 243180 68040 243306
rect 67158 242298 67284 243180
rect 67914 242298 68040 243180
rect 67158 242172 68040 242298
rect 65638 241794 67024 241920
rect 65638 241290 65764 241794
rect 66898 241290 67024 241794
rect 65638 241272 67024 241290
rect 65618 241112 67024 241272
rect 34295 240406 34647 240476
rect 34295 240344 34339 240406
rect 31908 239696 34339 240344
rect 34295 239180 34339 239696
rect 31908 238532 34339 239180
rect 7840 227920 20944 238448
rect 34295 237901 34339 238532
rect 31908 237262 34339 237901
rect 34594 237262 34647 240406
rect 31908 237253 34647 237262
rect 34295 237210 34647 237253
rect 67490 235372 67690 242172
rect 65347 235172 70972 235372
rect 65347 232265 65547 235172
rect 65347 232065 65547 232092
rect 65837 234573 68976 234773
rect 69088 234573 69129 234773
rect 65837 230800 66037 234573
rect 70772 234002 70972 235172
rect 66276 233604 66780 233730
rect 66276 232596 66402 233604
rect 66654 232596 66780 233604
rect 66276 232470 66780 232596
rect 65837 230600 66921 230800
rect 72324 229320 73710 229446
rect 66713 228483 66913 228926
rect 72324 228880 72450 229320
rect 69211 228483 69411 228840
rect 70732 228720 72450 228880
rect 72324 228690 72450 228720
rect 73584 228690 73710 229320
rect 72324 228564 73710 228690
rect 66713 228283 69411 228483
rect 493584 227136 506688 237664
rect 477520 225218 477548 225324
rect 477644 225218 477656 225324
rect 477712 225200 477862 225328
rect 477984 225200 478004 225328
rect 477982 224992 482160 225008
rect 477502 224880 477548 224992
rect 477644 224896 482160 224992
rect 482216 224896 482608 225008
rect 477644 224880 478114 224896
rect 477531 224274 477552 224396
rect 477648 224358 478114 224396
rect 477648 224274 478646 224358
rect 477989 224236 478646 224274
rect 478702 224236 482640 224358
rect 477538 223786 477552 223892
rect 477648 223786 477674 223892
rect 477736 223776 477862 223904
rect 477984 223776 478006 223904
rect 33126 223242 33425 223279
rect 31944 223223 33439 223242
rect 31944 222806 33176 223223
rect 33126 222454 33176 222806
rect 31954 222018 33176 222454
rect 7840 211120 20944 221648
rect 33126 220589 33176 222018
rect 31954 220153 33176 220589
rect 33126 219793 33176 220153
rect 31954 219357 33176 219793
rect 33382 222806 33439 223223
rect 33382 222454 33425 222806
rect 33382 222018 33439 222454
rect 33382 220589 33425 222018
rect 33382 220153 33439 220589
rect 33382 219793 33425 220153
rect 33382 219357 33439 219793
rect 33126 219314 33425 219357
rect 471904 211988 482633 212980
rect 471904 210668 482633 211660
rect 72828 209538 73710 209664
rect 72828 208656 72954 209538
rect 73584 208656 73710 209538
rect 471904 209348 482633 210340
rect 72828 208530 73710 208656
rect 72828 208476 73332 208530
rect 471904 208028 482633 209020
rect 79254 207942 79758 208026
rect 79254 207037 79331 207942
rect 79238 206980 79331 207037
rect 79685 207037 79758 207942
rect 79685 206980 79776 207037
rect 79238 206877 79776 206980
rect 34895 206806 35247 206876
rect 34895 206744 34939 206806
rect 31908 206096 34939 206744
rect 34895 205580 34939 206096
rect 31908 204932 34939 205580
rect 7840 194320 20944 204848
rect 34895 204301 34939 204932
rect 31908 203662 34939 204301
rect 35194 203662 35247 206806
rect 471904 206424 482633 207416
rect 74306 205722 74654 205762
rect 74306 205038 74345 205722
rect 74614 205038 74654 205722
rect 471904 205104 482633 206096
rect 74306 204864 74654 205038
rect 471904 203784 482633 204776
rect 31908 203653 35247 203662
rect 34895 203610 35247 203653
rect 471904 202180 482633 203172
rect 471904 200860 482633 201852
rect 471904 199540 482633 200532
rect 70686 198850 71442 198976
rect 70686 198094 70812 198850
rect 71316 198094 71442 198850
rect 471904 198220 482633 199212
rect 70686 197968 71442 198094
rect 68922 193032 69678 193158
rect 68922 192402 69048 193032
rect 69552 192402 69678 193032
rect 68922 192276 69678 192402
rect 69008 190924 69320 192276
rect 70898 191042 71098 197968
rect 471896 195188 482625 196180
rect 471896 193868 482625 194860
rect 471896 192548 482625 193540
rect 471896 191228 482625 192220
rect 35495 190006 35847 190076
rect 35495 189944 35539 190006
rect 31908 189296 35539 189944
rect 35495 188780 35539 189296
rect 31908 188132 35539 188780
rect 7840 177520 20944 188048
rect 35495 187501 35539 188132
rect 31908 186862 35539 187501
rect 35794 186862 35847 190006
rect 66024 190008 66906 190134
rect 66024 189252 66150 190008
rect 66780 189982 66906 190008
rect 66780 189252 67026 189982
rect 471896 189624 482625 190616
rect 66024 189140 67026 189252
rect 66024 189126 66906 189140
rect 471896 188304 482625 189296
rect 64473 187664 64545 187864
rect 64831 187664 67026 187864
rect 471896 186984 482625 187976
rect 31908 186853 35847 186862
rect 35495 186810 35847 186853
rect 66770 185968 67122 185991
rect 66770 185801 66801 185968
rect 67096 185801 67122 185968
rect 66770 185782 67122 185801
rect 471896 185380 482625 186372
rect 471896 184060 482625 185052
rect 471896 182740 482625 183732
rect 471896 181420 482625 182412
rect 36095 173206 36447 173276
rect 36095 173144 36139 173206
rect 31908 172496 36139 173144
rect 36095 171980 36139 172496
rect 31908 171332 36139 171980
rect 7840 160720 20944 171248
rect 36095 170701 36139 171332
rect 31908 170062 36139 170701
rect 36394 170062 36447 173206
rect 31908 170053 36447 170062
rect 36095 170010 36447 170053
rect 72828 167202 74214 167328
rect 72828 166446 73332 167202
rect 74088 166446 74214 167202
rect 72828 166320 74214 166446
rect 72828 166312 73332 166320
rect 79380 165312 80010 165438
rect 79380 164215 79506 165312
rect 79370 164178 79506 164215
rect 79884 164178 80010 165312
rect 79370 164055 80010 164178
rect 79380 164052 80010 164055
rect 80760 162040 81648 162200
rect 80766 162036 81648 162040
rect 80766 161532 80892 162036
rect 81522 161532 81648 162036
rect 80766 161406 81648 161532
rect 36695 156406 37047 156476
rect 36695 156344 36739 156406
rect 31935 155696 36739 156344
rect 36695 155180 36739 155696
rect 31944 154532 36739 155180
rect 7840 143920 20944 154448
rect 36695 153901 36739 154532
rect 31961 153262 36739 153901
rect 36994 153262 37047 156406
rect 31961 153253 37047 153262
rect 36695 153210 37047 153253
rect 51282 153468 52920 153594
rect 51282 152838 51408 153468
rect 52794 152838 52920 153468
rect 51282 152712 52920 152838
rect 51580 148712 51740 152712
rect 321000 149736 321600 149836
rect 321000 149336 321100 149736
rect 321500 149336 321600 149736
rect 321000 149236 321600 149336
rect 321100 148772 321500 149236
rect 51580 148552 52291 148712
rect 51580 146183 51740 148552
rect 52164 148371 52220 148385
rect 52164 148212 52220 148226
rect 52724 148370 52780 148384
rect 52724 148212 52780 148226
rect 53284 148370 53340 148384
rect 53284 148212 53340 148226
rect 53844 148370 53900 148384
rect 54188 147656 60560 147816
rect 60400 147079 60560 147656
rect 54054 146919 60560 147079
rect 52500 146848 52556 146861
rect 52500 146689 52556 146702
rect 53060 146848 53116 146861
rect 53060 146689 53116 146702
rect 53620 146848 53676 146861
rect 53620 146689 53676 146702
rect 54180 146848 54236 146861
rect 54180 146689 54236 146702
rect 50828 145568 51180 146024
rect 51580 146023 54270 146183
rect 60400 145404 60560 146919
rect 81144 146412 81774 146538
rect 60354 145400 60858 145404
rect 60354 145240 61488 145400
rect 60354 137088 60858 145240
rect 61684 145040 61740 145076
rect 61236 144890 61334 144966
rect 61390 144890 61404 144966
rect 61684 144773 61740 144816
rect 81144 144504 81270 146412
rect 79884 144344 81270 144504
rect 81144 142380 81270 144344
rect 81648 142380 81774 146412
rect 84818 145576 89792 145736
rect 84422 145361 84478 145412
rect 84422 145167 84478 145174
rect 86718 145202 86907 145353
rect 82432 144978 83216 145040
rect 82432 144633 82494 144978
rect 83152 144840 83216 144978
rect 83152 144680 86514 144840
rect 83152 144633 83216 144680
rect 82432 144592 83216 144633
rect 81144 142254 81774 142380
rect 89632 139440 89792 145576
rect 481824 144704 481908 144816
rect 481964 144704 482608 144816
rect 481824 144144 481908 144256
rect 481964 144144 482608 144256
rect 89152 139328 90832 139440
rect 89152 138432 89264 139328
rect 90720 138432 90832 139328
rect 480372 139324 480410 139446
rect 480466 139324 482640 139446
rect 89152 138320 90832 138432
rect 481824 138096 481908 138208
rect 481964 138096 482608 138208
rect 60354 136584 61488 137088
rect 493584 136752 506688 147280
rect 60858 135880 61488 136584
rect 81144 136458 81774 136584
rect 60858 135828 62118 135880
rect 60858 133560 60984 135828
rect 61362 135720 62118 135828
rect 61362 133640 61488 135720
rect 81144 134984 81270 136458
rect 79758 134946 81270 134984
rect 81648 134946 81774 136458
rect 481348 134952 481376 135058
rect 481472 134952 481484 135058
rect 79758 134824 81774 134946
rect 481540 134934 481690 135062
rect 481812 134934 481832 135062
rect 81144 134820 81774 134824
rect 479868 134444 479906 134566
rect 479962 134444 481376 134566
rect 481472 134444 482640 134566
rect 480120 133956 480158 134078
rect 480214 133956 481380 134078
rect 481476 133956 482640 134078
rect 275800 133700 276600 133800
rect 61362 133560 61822 133640
rect 60858 133480 61822 133560
rect 60858 133434 61488 133480
rect 61030 131287 61190 133434
rect 275800 133100 275900 133700
rect 276500 133100 276600 133700
rect 481366 133520 481380 133626
rect 481476 133520 481502 133626
rect 481564 133510 481690 133638
rect 481812 133510 481834 133638
rect 275800 133000 276600 133100
rect 72188 132804 73196 132930
rect 72188 132744 72314 132804
rect 66448 132584 72314 132744
rect 72188 132174 72314 132584
rect 73070 132174 73196 132804
rect 276000 132200 276400 133000
rect 72188 132048 73196 132174
rect 62622 131292 65772 131418
rect 62622 131287 62748 131292
rect 60400 131127 62748 131287
rect 62622 131040 62748 131127
rect 65646 131040 65772 131292
rect 62622 130914 65772 131040
rect 62622 130410 65772 130536
rect 62622 130391 62748 130410
rect 61962 130390 62748 130391
rect 61874 130231 62748 130390
rect 62622 130158 62748 130231
rect 65646 130158 65772 130410
rect 62622 130032 65772 130158
rect 481824 127904 481908 128016
rect 481964 127904 482608 128016
rect 7840 117152 20944 127680
rect 59724 127652 60228 127764
rect 59014 127638 60228 127652
rect 59014 127492 59850 127638
rect 59724 127386 59850 127492
rect 60102 127386 60228 127638
rect 59724 127260 60228 127386
rect 481824 127344 481908 127456
rect 481964 127344 482608 127456
rect 59101 127246 59243 127247
rect 59101 127082 59115 127246
rect 59193 127082 59243 127246
rect 60984 127008 61992 127134
rect 60984 126676 61110 127008
rect 59012 126630 61110 126676
rect 61866 126630 61992 127008
rect 117420 126788 117460 126844
rect 117516 126788 119952 126844
rect 59012 126516 61992 126630
rect 60984 126504 61992 126516
rect 117644 125780 117684 125836
rect 117740 125780 119979 125836
rect 479112 122488 479150 122610
rect 479206 122488 482640 122610
rect 481824 121296 481908 121408
rect 481964 121296 482608 121408
rect 493584 119952 506688 130480
rect 117868 119844 117908 119900
rect 117964 119844 119979 119900
rect 118092 118948 118132 119004
rect 118188 118948 119979 119004
rect 481348 118152 481376 118258
rect 481472 118152 481484 118258
rect 481540 118134 481690 118262
rect 481812 118134 481832 118262
rect 118316 117940 118356 117996
rect 118412 117940 119979 117996
rect 479616 117730 479654 117852
rect 479710 117730 481376 117852
rect 481472 117730 482640 117852
rect 479364 117120 479402 117242
rect 479458 117120 481380 117242
rect 481476 117120 482640 117242
rect 118540 116932 118580 116988
rect 118636 116932 119979 116988
rect 481366 116720 481380 116826
rect 481476 116720 481502 116826
rect 481564 116710 481690 116838
rect 481812 116710 481834 116838
rect 31962 115067 112015 115954
rect 118764 115924 118804 115980
rect 118860 115924 119979 115980
rect 69634 111844 72178 112004
rect 71972 111820 72178 111844
rect 37548 109620 39186 109746
rect 37548 108612 37674 109620
rect 38556 108612 39186 109620
rect 66740 109242 67340 111022
rect 71972 109531 72179 111820
rect 89694 110100 92584 110300
rect 91302 109620 91902 109794
rect 37548 108486 39186 108612
rect 60022 109056 64263 109216
rect 66740 109116 67662 109242
rect 71972 109224 74940 109531
rect 91302 109418 91476 109620
rect 60022 108974 62110 109056
rect 38504 105966 39104 108486
rect 60022 107478 60182 108974
rect 66740 108738 66906 109116
rect 67536 108738 67662 109116
rect 70858 109064 74940 109224
rect 89690 109218 91476 109418
rect 66740 108612 67662 108738
rect 61972 108534 63460 108590
rect 66740 108248 67340 108612
rect 68135 108469 68152 108581
rect 68212 108469 68232 108581
rect 68903 108527 69183 108621
rect 61416 108088 71648 108248
rect 65772 107604 66680 107730
rect 59472 107352 60732 107478
rect 59472 106974 59598 107352
rect 60606 106974 60732 107352
rect 65772 107226 65898 107604
rect 66528 107226 66680 107604
rect 65772 107100 66680 107226
rect 59472 106848 60732 106974
rect 59760 105966 60360 106848
rect 66080 105966 66680 107100
rect 66740 105966 67340 108088
rect 74505 107982 74940 109064
rect 86397 108538 86412 108738
rect 86640 108538 86888 108738
rect 89707 108424 89839 109218
rect 91302 108738 91476 109218
rect 91728 108738 91902 109620
rect 74214 107856 75222 107982
rect 74214 107352 74340 107856
rect 75096 107352 75222 107856
rect 90342 107856 90972 107982
rect 90342 107608 90468 107856
rect 89698 107478 90468 107608
rect 90846 107478 90972 107856
rect 89698 107408 90972 107478
rect 90342 107352 90972 107408
rect 74214 107226 75222 107352
rect 74074 107072 74196 107086
rect 74074 105963 74196 107016
rect 74416 105966 75016 107226
rect 91302 107100 91902 108738
rect 92384 107982 92584 110100
rect 92358 107856 93114 107982
rect 92358 107352 92484 107856
rect 92988 107352 93114 107856
rect 92358 107226 93114 107352
rect 89730 106422 91902 107100
rect 89730 105966 90330 106422
rect 31708 95508 35188 95584
rect 35244 95508 35284 95584
rect 31708 78102 35524 78178
rect 35580 78102 35616 78178
rect 111128 74276 112015 115067
rect 118988 114916 119028 114972
rect 119084 114916 119979 114972
rect 116524 114020 116564 114076
rect 116620 114020 119979 114076
rect 116300 113012 116340 113068
rect 116396 113012 119979 113068
rect 117196 112004 117236 112060
rect 117292 112004 119979 112060
rect 117420 111444 117460 111500
rect 117516 111444 119979 111500
rect 117644 109988 117684 110044
rect 117740 109988 119979 110044
rect 117868 108448 117908 108504
rect 117964 108448 119979 108504
rect 118092 106992 118132 107048
rect 118188 106992 119979 107048
rect 477300 78500 477700 78974
rect 477200 78400 477800 78500
rect 477200 78000 477300 78400
rect 477700 78000 477800 78400
rect 477200 77900 477800 78000
rect 472400 75780 478000 75800
rect 472400 75600 482618 75780
rect 111128 73389 198741 74276
rect 119236 72760 119264 72820
rect 119904 72760 120274 72820
rect 119244 72600 119264 72660
rect 119904 72600 120274 72660
rect 114597 72198 115227 72261
rect 113148 72072 114030 72198
rect 113148 71442 113274 72072
rect 113904 71442 114030 72072
rect 114597 71694 114660 72198
rect 115164 72168 115227 72198
rect 115164 72070 120526 72168
rect 115164 72008 120686 72070
rect 133300 72828 140986 72954
rect 115164 71694 115227 72008
rect 114597 71631 115227 71694
rect 116056 71564 116067 71620
rect 116239 71564 116250 71620
rect 133300 71442 136072 72828
rect 140860 71442 140986 72828
rect 113148 71318 116046 71442
rect 113148 71316 114030 71318
rect 133300 71316 140986 71442
rect 133300 71272 134938 71316
rect 117226 71112 134938 71272
rect 133300 70560 134938 71112
rect 133472 70480 133632 70560
rect 197854 59885 198741 73389
rect 268380 61362 283248 61488
rect 197854 59840 206712 59885
rect 197854 59033 205006 59840
rect 206669 59033 206712 59840
rect 268380 59472 268506 61362
rect 283122 59472 283248 61362
rect 472400 61200 472600 75600
rect 477800 74788 482618 75600
rect 477800 74460 478000 74788
rect 477800 73468 482618 74460
rect 477800 73140 478000 73468
rect 477800 72148 482618 73140
rect 477800 71820 478000 72148
rect 477800 70828 482618 71820
rect 477800 70216 478000 70828
rect 477800 69224 482618 70216
rect 477800 68896 478000 69224
rect 477800 67904 482618 68896
rect 477800 67576 478000 67904
rect 477800 66584 482618 67576
rect 477800 65972 478000 66584
rect 477800 64980 482618 65972
rect 477800 64652 478000 64980
rect 477800 63660 482618 64652
rect 477800 63332 478000 63660
rect 477800 62340 482618 63332
rect 477800 62012 478000 62340
rect 477800 61200 482618 62012
rect 472400 61020 482618 61200
rect 472400 61000 478000 61020
rect 268380 59346 283248 59472
rect 197854 58998 206712 59033
rect 34400 57780 36400 57800
rect 31947 57600 36400 57780
rect 31947 56788 34600 57600
rect 34400 56460 34600 56788
rect 31947 55468 34600 56460
rect 34400 55140 34600 55468
rect 31947 54148 34600 55140
rect 34400 53820 34600 54148
rect 31947 52828 34600 53820
rect 34400 52216 34600 52828
rect 31947 51224 34600 52216
rect 34400 50896 34600 51224
rect 31947 49904 34600 50896
rect 34400 49576 34600 49904
rect 31947 48584 34600 49576
rect 34400 47972 34600 48584
rect 31947 46980 34600 47972
rect 34400 46652 34600 46980
rect 31947 45660 34600 46652
rect 34400 45332 34600 45660
rect 31947 44340 34600 45332
rect 34400 44012 34600 44340
rect 31947 43200 34600 44012
rect 36200 43200 36400 57600
rect 199000 53800 204646 54000
rect 199000 51600 199200 53800
rect 204464 51600 204646 53800
rect 199000 51400 204646 51600
rect 199052 51322 204646 51400
rect 205266 53800 211000 54000
rect 205266 51600 205440 53800
rect 210800 51600 211000 53800
rect 205266 51400 211000 51600
rect 205266 51322 210864 51400
rect 199052 50633 204652 51322
rect 205264 50633 210864 51322
rect 31947 43020 36400 43200
rect 34400 43000 36400 43020
rect 231600 42200 246400 42400
rect 59700 41700 60500 41800
rect 59700 41100 59800 41700
rect 60400 41100 60500 41700
rect 59700 41000 60500 41100
rect 59900 40464 60300 41000
rect 231600 37200 231800 42200
rect 246200 37200 246400 42200
rect 231600 37000 246400 37200
rect 102200 35400 117000 35600
rect 34992 34184 35048 34254
rect 34362 33932 34418 33944
rect 34362 31936 34418 33876
rect 34992 31936 35048 34128
rect 102200 33800 102400 35400
rect 116800 33800 117000 35400
rect 73422 33680 73478 33720
rect 56538 33428 56594 33468
rect 55404 32680 55460 32720
rect 55404 31936 55460 32624
rect 56538 31936 56594 33372
rect 72162 32680 72218 32720
rect 72162 31936 72218 32624
rect 73422 31936 73478 33624
rect 102200 33600 117000 33800
rect 90180 33176 90236 33216
rect 88920 32680 88976 32720
rect 88920 31936 88976 32624
rect 90180 31936 90236 33120
rect 102220 31952 103212 33600
rect 103540 31952 104532 33600
rect 104860 31952 105852 33600
rect 106180 31952 107172 33600
rect 107784 31952 108776 33600
rect 109104 31952 110096 33600
rect 110424 31952 111416 33600
rect 112028 31952 113020 33600
rect 113348 31952 114340 33600
rect 114668 31952 115660 33600
rect 115988 31952 116980 33600
rect 231620 31920 232612 37000
rect 232940 31920 233932 37000
rect 234260 31920 235252 37000
rect 235580 31920 236572 37000
rect 237184 31920 238176 37000
rect 238504 31920 239496 37000
rect 239824 31920 240816 37000
rect 241428 31920 242420 37000
rect 242748 31920 243740 37000
rect 244068 31920 245060 37000
rect 245388 31920 246380 37000
rect 268420 31962 269412 59346
rect 269740 31962 270732 59346
rect 271060 31962 272052 59346
rect 272380 31962 273372 59346
rect 273984 31962 274976 59346
rect 275304 31962 276296 59346
rect 276624 31962 277616 59346
rect 278228 31962 279220 59346
rect 279548 31962 280540 59346
rect 280868 31962 281860 59346
rect 282188 31962 283180 59346
rect 285200 58600 300000 58800
rect 285200 53400 285400 58600
rect 299800 53400 300000 58600
rect 285200 53200 300000 53400
rect 285220 31939 286212 53200
rect 286540 31939 287532 53200
rect 287860 31939 288852 53200
rect 289180 31939 290172 53200
rect 290784 31939 291776 53200
rect 292104 31939 293096 53200
rect 293424 31939 294416 53200
rect 295028 31939 296020 53200
rect 296348 31939 297340 53200
rect 297668 31939 298660 53200
rect 298988 31939 299980 53200
rect 318000 51200 318400 51762
rect 317800 51100 318600 51200
rect 317800 50500 317900 51100
rect 318500 50500 318600 51100
rect 317800 50400 318600 50500
rect 481320 48922 481418 49044
rect 481474 48922 482640 49044
rect 481824 47712 481908 47824
rect 481964 47712 482608 47824
rect 493584 46368 506688 56896
rect 480596 43800 481018 44577
rect 480400 43700 481200 43800
rect 480400 43100 480500 43700
rect 481100 43100 481200 43700
rect 480400 43000 481200 43100
rect 328104 37604 328230 37698
rect 311346 36384 311472 36478
rect 310886 33200 311014 33222
rect 310886 32952 311014 33078
rect 310896 32864 311002 32890
rect 310896 32754 311002 32768
rect 311346 32864 311472 36328
rect 311346 31964 311472 32768
rect 311976 36140 312102 36234
rect 311976 32860 312102 36084
rect 312310 33200 312438 33220
rect 312310 32928 312438 33078
rect 327686 33200 327814 33222
rect 327686 32952 327814 33078
rect 311976 31964 312102 32764
rect 312328 32860 312434 32872
rect 312328 32736 312434 32764
rect 327696 32864 327802 32890
rect 327696 32754 327802 32768
rect 328104 32864 328230 37548
rect 420714 37360 420840 37454
rect 403956 37116 404082 37210
rect 387072 36872 387198 36966
rect 370314 36628 370440 36722
rect 328104 31964 328230 32768
rect 328734 35896 328860 35990
rect 328734 32860 328860 35840
rect 365526 35652 365652 35746
rect 364896 34686 365022 34770
rect 329110 33200 329238 33220
rect 329110 32928 329238 33078
rect 364486 33200 364614 33222
rect 364486 32952 364614 33078
rect 328734 31964 328860 32764
rect 329128 32860 329234 32872
rect 329128 32736 329234 32764
rect 364496 32864 364602 32890
rect 364496 32754 364602 32768
rect 364896 32864 365022 34630
rect 364896 31964 365022 32768
rect 365526 32860 365652 35596
rect 369040 33404 369152 33488
rect 365910 33200 366038 33220
rect 365910 32928 366038 33078
rect 365526 31964 365652 32764
rect 365928 32860 366034 32872
rect 365928 32736 366034 32764
rect 369040 31920 369152 33348
rect 370314 31964 370440 36572
rect 382284 35408 382410 35502
rect 381654 34434 381780 34526
rect 381286 33200 381414 33222
rect 381286 32952 381414 33078
rect 381296 32864 381402 32890
rect 381296 32754 381402 32768
rect 381654 32864 381780 34378
rect 381654 31964 381780 32768
rect 382284 32860 382410 35352
rect 385840 33404 385952 33488
rect 382710 33200 382838 33220
rect 382710 32928 382838 33078
rect 382284 31964 382410 32764
rect 382728 32860 382834 32872
rect 382728 32736 382834 32764
rect 385840 31920 385952 33348
rect 387072 31964 387198 36816
rect 399168 35164 399294 35258
rect 398538 34182 398664 34282
rect 398086 33200 398214 33222
rect 398086 32952 398214 33078
rect 398096 32864 398202 32890
rect 398096 32754 398202 32768
rect 398538 32864 398664 34126
rect 398538 31964 398664 32768
rect 399168 32860 399294 35108
rect 402640 33404 402752 33488
rect 399510 33200 399638 33220
rect 399510 32928 399638 33078
rect 399168 31964 399294 32764
rect 399528 32860 399634 32872
rect 399528 32736 399634 32764
rect 402640 31920 402752 33348
rect 403956 31964 404082 37060
rect 415926 34980 416052 35074
rect 415296 33930 415422 34038
rect 414886 33200 415014 33222
rect 414886 32952 415014 33078
rect 414896 32864 415002 32890
rect 414896 32754 415002 32768
rect 415296 32864 415422 33874
rect 415296 31964 415422 32768
rect 415926 32860 416052 34924
rect 419440 33404 419552 33488
rect 416310 33200 416438 33220
rect 416310 32928 416438 33078
rect 415926 31964 416052 32764
rect 416328 32860 416434 32872
rect 416328 32736 416434 32764
rect 419440 31920 419552 33348
rect 420714 31964 420840 37304
rect 432820 33200 433812 38934
rect 432820 31922 433812 33078
rect 434140 31922 435132 38934
rect 435460 31922 436452 38934
rect 436780 31922 437772 38934
rect 438384 31922 439376 38934
rect 439704 31922 440696 38934
rect 441024 31922 442016 38934
rect 442628 31922 443620 38934
rect 443948 31922 444940 38934
rect 445268 31922 446260 38934
rect 446588 31922 447580 38934
rect 471492 33662 471618 33672
rect 470288 33404 470400 33488
rect 470288 31920 470400 33348
rect 471492 31964 471618 33606
rect 37136 7840 47664 20944
rect 53936 7840 64464 20944
rect 70736 7840 81264 20944
rect 87536 7840 98064 20944
rect 287280 7840 297808 20944
rect 314160 7840 324688 20944
rect 330960 7840 341488 20944
rect 367696 7840 378224 20944
rect 384496 7840 395024 20944
rect 401296 7840 411824 20944
rect 418096 7840 428624 20944
rect 468944 7840 479472 20944
<< via1 >>
rect 37520 380996 37632 381052
rect 33600 366000 34600 380400
rect 37070 378594 37160 378686
rect 37520 378594 37632 378686
rect 35550 378058 35872 378202
rect 38192 381108 38304 381164
rect 44128 381332 44240 381388
rect 43008 380772 43120 380828
rect 47712 380884 47824 380940
rect 38192 378568 38304 378660
rect 38666 378568 38756 378660
rect 47262 378594 47352 378686
rect 47712 378594 47824 378686
rect 48384 381220 48496 381276
rect 54320 380436 54432 380492
rect 48384 378568 48496 378660
rect 48858 378568 48948 378660
rect 53870 378594 53960 378686
rect 54320 378594 54432 378686
rect 54992 380548 55104 380604
rect 60928 381332 61040 381388
rect 59808 380212 59920 380268
rect 64512 380324 64624 380380
rect 54992 378568 55104 378660
rect 37050 378058 37182 378202
rect 38640 378058 38772 378202
rect 55466 378568 55556 378660
rect 64062 378594 64152 378686
rect 64512 378594 64624 378686
rect 65184 380660 65296 380716
rect 71120 379876 71232 379932
rect 65184 378568 65296 378660
rect 47242 378058 47374 378202
rect 48832 378058 48964 378202
rect 53850 378058 53982 378202
rect 55440 378058 55572 378202
rect 65658 378568 65748 378660
rect 70670 378594 70760 378686
rect 71120 378594 71232 378686
rect 71792 379988 71904 380044
rect 77728 381332 77840 381388
rect 76608 379652 76720 379708
rect 77110 380100 77228 380156
rect 71792 378568 71904 378660
rect 72266 378568 72356 378660
rect 76662 378594 76752 378686
rect 77112 378594 77224 378686
rect 77784 379764 77898 379820
rect 87470 380994 87560 381086
rect 87920 380994 88032 381086
rect 87450 380458 87582 380602
rect 81984 380100 82096 380156
rect 81312 379764 81424 379820
rect 88592 380968 88704 381060
rect 89066 380968 89156 381060
rect 89040 380458 89172 380602
rect 88592 379428 88704 379484
rect 87920 379316 88032 379372
rect 77784 378568 77896 378660
rect 78258 378568 78348 378660
rect 64042 378058 64174 378202
rect 65632 378058 65764 378202
rect 70650 378058 70782 378202
rect 72240 378058 72372 378202
rect 76642 378058 76774 378202
rect 78232 378058 78364 378202
rect 94528 381332 94640 381388
rect 97662 380994 97752 381086
rect 98112 380994 98224 381086
rect 97642 380458 97774 380602
rect 98784 380968 98896 381060
rect 99258 380968 99348 381060
rect 104270 380994 104360 381086
rect 104720 380994 104832 381086
rect 99232 380458 99364 380602
rect 104250 380458 104382 380602
rect 98784 379540 98896 379596
rect 98112 379204 98224 379260
rect 105392 380968 105504 381060
rect 105866 380968 105956 381060
rect 105840 380458 105972 380602
rect 105392 378980 105504 379036
rect 104720 378868 104832 378924
rect 93380 374257 93436 374927
rect 111328 381332 111440 381388
rect 114462 380994 114552 381086
rect 114912 380994 115024 381086
rect 114442 380458 114574 380602
rect 115584 380968 115696 381060
rect 116058 380968 116148 381060
rect 121070 380994 121160 381086
rect 121520 380994 121632 381086
rect 116032 380458 116164 380602
rect 121050 380458 121182 380602
rect 115584 379092 115696 379148
rect 114912 378756 115024 378812
rect 122192 380968 122304 381060
rect 122666 380968 122756 381060
rect 122640 380458 122772 380602
rect 122192 378532 122304 378588
rect 121520 378420 121632 378476
rect 110180 374257 110236 374927
rect 128128 381332 128240 381388
rect 131262 380994 131352 381086
rect 131712 380994 131824 381086
rect 131242 380458 131374 380602
rect 132384 380968 132496 381060
rect 132858 380968 132948 381060
rect 137870 380994 137960 381086
rect 138320 380994 138432 381086
rect 132832 380458 132964 380602
rect 137850 380458 137982 380602
rect 132384 378644 132496 378700
rect 131712 378308 131824 378364
rect 138992 380968 139104 381060
rect 139466 380968 139556 381060
rect 139440 380458 139572 380602
rect 138992 378084 139104 378140
rect 138320 377972 138432 378028
rect 126980 374257 127036 374927
rect 144928 381332 145040 381388
rect 148062 380994 148152 381086
rect 148512 380994 148624 381086
rect 148042 380458 148174 380602
rect 149184 380968 149296 381060
rect 149658 380968 149748 381060
rect 194670 380994 194760 381086
rect 195120 380994 195232 381086
rect 149632 380458 149764 380602
rect 194650 380458 194782 380602
rect 149184 378196 149296 378252
rect 148512 377860 148624 377916
rect 195792 380968 195904 381060
rect 196266 380968 196356 381060
rect 196240 380458 196372 380602
rect 195792 377636 195904 377692
rect 195120 377524 195232 377580
rect 143780 374257 143836 374927
rect 201712 381332 201824 381388
rect 204862 380994 204952 381086
rect 205312 380994 205424 381086
rect 204842 380458 204974 380602
rect 205984 380968 206096 381060
rect 206458 380968 206548 381060
rect 211470 380994 211560 381086
rect 211920 380994 212032 381086
rect 206432 380458 206564 380602
rect 211450 380458 211582 380602
rect 205984 377748 206096 377804
rect 205312 377412 205424 377468
rect 212592 380968 212704 381060
rect 213066 380968 213156 381060
rect 213040 380458 213172 380602
rect 212592 377188 212704 377244
rect 211920 377076 212032 377132
rect 200580 374257 200636 374927
rect 218512 381332 218624 381388
rect 221662 380994 221752 381086
rect 222112 380994 222224 381086
rect 221642 380458 221774 380602
rect 222784 380968 222896 381060
rect 223258 380968 223348 381060
rect 238270 380994 238360 381086
rect 238720 380994 238832 381086
rect 223232 380458 223364 380602
rect 238250 380458 238382 380602
rect 222784 377300 222896 377356
rect 222112 376964 222224 377020
rect 239392 380968 239504 381060
rect 239866 380968 239956 381060
rect 239840 380458 239972 380602
rect 239392 376740 239504 376796
rect 238720 376628 238832 376684
rect 217380 374257 217436 374927
rect 245280 381332 245392 381388
rect 248462 380994 248552 381086
rect 248912 380994 249024 381086
rect 248442 380458 248574 380602
rect 249584 380968 249696 381060
rect 250058 380968 250148 381060
rect 255070 380994 255160 381086
rect 255520 380994 255632 381086
rect 250032 380458 250164 380602
rect 255050 380458 255182 380602
rect 249584 376852 249696 376908
rect 248912 376516 249024 376572
rect 256192 380968 256304 381060
rect 256666 380968 256756 381060
rect 256640 380458 256772 380602
rect 256192 376292 256304 376348
rect 255520 376180 255632 376236
rect 244180 374257 244236 374927
rect 262080 381332 262192 381388
rect 265262 380994 265352 381086
rect 265712 380994 265824 381086
rect 265242 380458 265374 380602
rect 266384 380968 266496 381060
rect 266858 380968 266948 381060
rect 271870 380994 271960 381086
rect 272320 380994 272432 381086
rect 266832 380458 266964 380602
rect 271850 380458 271982 380602
rect 266384 376404 266496 376460
rect 265712 376068 265824 376124
rect 272992 380968 273104 381060
rect 273466 380968 273556 381060
rect 273440 380458 273572 380602
rect 272992 375844 273104 375900
rect 272320 375732 272432 375788
rect 260980 374257 261036 374927
rect 278880 381332 278992 381388
rect 282062 380994 282152 381086
rect 282512 380994 282624 381086
rect 282042 380458 282174 380602
rect 283184 380968 283296 381060
rect 283658 380968 283748 381060
rect 283632 380458 283764 380602
rect 283184 375956 283296 376012
rect 282512 375620 282624 375676
rect 277780 374257 277836 374927
rect 427400 374200 441800 375800
rect 444200 374200 458600 375800
rect 467000 374200 481400 375800
rect 470383 373083 470645 373345
rect 471500 373000 472000 373500
rect 480662 370514 480718 370636
rect 481908 369264 481964 369376
rect 33600 349200 34600 363600
rect 63504 366912 64764 367542
rect 320796 364604 322686 365486
rect 328783 364983 329045 365245
rect 328600 363400 329200 364000
rect 65394 360360 65646 360864
rect 66150 360360 66780 361620
rect 320684 362847 320740 363034
rect 321020 362908 321188 362964
rect 322056 361872 323316 362502
rect 319645 361252 319701 361422
rect 321040 361265 321096 361525
rect 316890 360612 317646 360990
rect 334600 360800 346000 362200
rect 63478 359934 63542 360122
rect 64778 360116 64940 360172
rect 63126 358092 63378 358470
rect 63662 358418 63798 358494
rect 64092 358367 64148 358554
rect 64332 358418 64472 358494
rect 64764 358367 64820 358554
rect 272636 357390 272692 357648
rect 272888 357390 272944 357648
rect 273140 357390 273196 357648
rect 273392 357390 273448 357648
rect 273644 357390 273700 357648
rect 273896 357390 273952 357648
rect 274148 357390 274204 357648
rect 89824 356090 90170 356146
rect 89824 355846 90170 355902
rect 89824 355602 90170 355658
rect 89824 355358 90170 355414
rect 89824 355114 90170 355170
rect 89824 354870 90170 354926
rect 89824 354626 90170 354682
rect 89824 354382 90170 354438
rect 89824 354138 90170 354194
rect 89824 353894 90170 353950
rect 472600 349200 477800 363600
rect 410256 340578 411894 341712
rect 32808 338042 32900 338132
rect 33226 338016 33370 338148
rect 32808 337568 32900 337680
rect 34020 337568 34076 337680
rect 32782 337008 32874 337120
rect 34356 337008 34412 337120
rect 32782 336558 32874 336648
rect 33226 336538 33370 336670
rect 32228 333312 32284 333424
rect 477548 332418 477644 332524
rect 477862 332400 477984 332528
rect 34468 332192 34524 332304
rect 477548 332080 477644 332192
rect 482160 332080 482216 332192
rect 477552 331474 477648 331596
rect 481166 331474 481222 331596
rect 477552 330986 477648 331092
rect 477862 330976 477984 331104
rect 32808 327850 32900 327940
rect 33226 327824 33370 327956
rect 32808 327376 32900 327488
rect 34132 327376 34188 327488
rect 32782 326704 32874 326816
rect 34244 326704 34300 326816
rect 32782 326254 32874 326344
rect 33226 326234 33370 326366
rect 32808 321242 32900 321332
rect 33226 321216 33370 321348
rect 32808 320768 32900 320880
rect 33460 320768 33516 320880
rect 32782 320208 32874 320320
rect 33796 320208 33852 320320
rect 32782 319758 32874 319848
rect 33226 319738 33370 319870
rect 332990 316684 333046 316862
rect 32228 316512 32284 316624
rect 333368 316684 333424 316862
rect 333872 316684 333928 316862
rect 336644 316684 336700 316862
rect 337148 316684 337204 316862
rect 337652 316684 337708 316862
rect 340424 316684 340480 316862
rect 340928 316684 340984 316862
rect 341432 316684 341488 316862
rect 344204 316684 344260 316862
rect 344708 316684 344764 316862
rect 345212 316684 345268 316862
rect 347984 316684 348040 316862
rect 348488 316684 348544 316862
rect 348992 316684 349048 316862
rect 351764 316684 351820 316862
rect 352268 316684 352324 316862
rect 352772 316684 352828 316862
rect 355544 316684 355600 316862
rect 356048 316684 356104 316862
rect 356552 316684 356608 316862
rect 359324 316684 359380 316862
rect 359828 316684 359884 316862
rect 360332 316684 360388 316862
rect 363104 316684 363160 316862
rect 363608 316684 363664 316862
rect 364112 316684 364168 316862
rect 366758 316684 366814 316862
rect 367262 316684 367318 316862
rect 367766 316684 367822 316862
rect 370538 316684 370594 316862
rect 371042 316684 371098 316862
rect 371546 316684 371602 316862
rect 374318 316684 374374 316862
rect 374822 316684 374878 316862
rect 375326 316684 375382 316862
rect 378098 316684 378154 316862
rect 378602 316684 378658 316862
rect 379106 316684 379162 316862
rect 381878 316684 381934 316862
rect 382382 316684 382438 316862
rect 382886 316684 382942 316862
rect 385658 316684 385714 316862
rect 386162 316684 386218 316862
rect 386666 316684 386722 316862
rect 389438 316684 389494 316862
rect 389942 316684 389998 316862
rect 390446 316684 390502 316862
rect 395612 316684 395668 316862
rect 396116 316684 396172 316862
rect 396872 316684 396928 316862
rect 398006 316684 398062 316862
rect 401534 316684 401590 316862
rect 402038 316684 402094 316862
rect 402542 316684 402598 316862
rect 403046 316684 403102 316862
rect 403550 316684 403606 316862
rect 404054 316684 404110 316862
rect 404558 316684 404614 316862
rect 405062 316684 405118 316862
rect 405566 316684 405622 316862
rect 406070 316684 406126 316862
rect 408842 316684 408898 316862
rect 409346 316684 409402 316862
rect 409850 316684 409906 316862
rect 412622 316684 412678 316862
rect 413126 316684 413182 316862
rect 413630 316684 413686 316862
rect 416402 316684 416458 316862
rect 416906 316684 416962 316862
rect 417410 316684 417466 316862
rect 420182 316684 420238 316862
rect 420686 316684 420742 316862
rect 421190 316684 421246 316862
rect 423962 316684 424018 316862
rect 424466 316684 424522 316862
rect 424970 316684 425026 316862
rect 427616 316684 427672 316862
rect 428120 316684 428176 316862
rect 428624 316684 428680 316862
rect 431396 316684 431452 316862
rect 431900 316684 431956 316862
rect 432404 316684 432460 316862
rect 435176 316684 435232 316862
rect 435680 316684 435736 316862
rect 436184 316684 436240 316862
rect 438956 316684 439012 316862
rect 439460 316684 439516 316862
rect 439964 316684 440020 316862
rect 442736 316684 442792 316862
rect 443240 316684 443296 316862
rect 443744 316684 443800 316862
rect 446516 316684 446572 316862
rect 447020 316684 447076 316862
rect 447524 316684 447580 316862
rect 450296 316684 450352 316862
rect 450800 316684 450856 316862
rect 451304 316684 451360 316862
rect 454076 316684 454132 316862
rect 454580 316684 454636 316862
rect 455084 316684 455140 316862
rect 457730 316684 457786 316862
rect 458234 316684 458290 316862
rect 458738 316684 458794 316862
rect 461510 316684 461566 316862
rect 462014 316684 462070 316862
rect 462518 316684 462574 316862
rect 465290 316684 465346 316862
rect 465794 316684 465850 316862
rect 466298 316684 466354 316862
rect 477548 315618 477644 315724
rect 477862 315600 477984 315728
rect 33908 315392 33964 315504
rect 477548 315280 477644 315392
rect 482160 315280 482216 315392
rect 477552 314674 477648 314796
rect 481418 314760 481474 314882
rect 477552 314186 477648 314292
rect 477862 314176 477984 314304
rect 35154 312984 35910 313488
rect 38413 313438 38578 313604
rect 39889 313438 40051 313597
rect 41744 313438 41962 313623
rect 42840 312858 43218 313614
rect 45467 313456 45631 313601
rect 46935 313456 47111 313610
rect 48779 313456 49011 313634
rect 60354 313110 61236 313362
rect 62636 312956 62804 313012
rect 63084 312886 63140 313073
rect 64512 312480 65394 312732
rect 32808 311050 32900 311140
rect 33226 311024 33370 311156
rect 32808 310576 32900 310688
rect 33572 310576 33628 310688
rect 42840 310338 43218 310842
rect 50022 310338 50400 310842
rect 32782 309904 32874 310016
rect 33684 309904 33740 310016
rect 32782 309454 32874 309544
rect 33226 309434 33370 309566
rect 60354 311220 61236 311850
rect 62734 311337 62798 311525
rect 64135 311287 64192 311457
rect 64526 311307 64590 311555
rect 65927 311287 65984 311457
rect 66320 311445 66380 311576
rect 67719 311287 67776 311457
rect 64184 311041 64240 311165
rect 65976 311041 66032 311165
rect 67768 311041 67824 311165
rect 68670 310968 69426 311220
rect 52708 310398 52947 310598
rect 50652 309078 51282 309582
rect 57903 310206 58105 310424
rect 68976 310214 69088 310414
rect 58590 308952 58842 309582
rect 53900 308460 54100 308560
rect 32358 304430 32430 304556
rect 32566 304462 32632 304526
rect 32566 303968 32632 304080
rect 32900 303968 32956 304080
rect 32540 303408 32612 303520
rect 33236 303408 33292 303520
rect 32358 302836 32438 302962
rect 32540 302860 32612 302936
rect 32228 299712 32284 299824
rect 477548 298818 477644 298924
rect 477862 298800 477984 298928
rect 33348 298592 33404 298704
rect 477548 298480 477644 298592
rect 481670 298534 481726 298656
rect 477552 297874 477648 297996
rect 480914 297924 480970 298046
rect 477552 297386 477648 297492
rect 477862 297376 477984 297504
rect 32358 294118 32448 294244
rect 32562 294140 32630 294224
rect 32562 293776 32630 293888
rect 33012 293776 33068 293888
rect 32540 293104 32610 293216
rect 33124 293104 33180 293216
rect 32358 292524 32434 292650
rect 32540 292546 32610 292630
rect 32358 288570 32454 288694
rect 32570 288596 32656 288670
rect 32108 288270 32164 288326
rect 32570 288270 32656 288326
rect 32358 287776 32446 287904
rect 32554 287804 32628 287882
rect 32108 287168 32164 287280
rect 32340 287168 32396 287280
rect 32554 286608 32628 286720
rect 32676 286608 32732 286720
rect 32228 282912 32284 283024
rect 32788 281792 32844 281904
rect 33108 277450 33200 277540
rect 33526 277424 33670 277556
rect 32452 276976 32508 277088
rect 33108 276976 33200 277088
rect 32564 276304 32620 276416
rect 33082 276304 33174 276416
rect 33082 275854 33174 275944
rect 33526 275834 33670 275966
rect 33739 254062 33994 257206
rect 478898 246440 478954 246562
rect 481908 245280 481964 245392
rect 63882 243936 64638 244692
rect 67284 242298 67914 243180
rect 65764 241290 66898 241794
rect 34339 237262 34594 240406
rect 65347 232092 65547 232265
rect 68976 234573 69088 234773
rect 66402 232596 66654 233604
rect 72450 228690 73584 229320
rect 477548 225218 477644 225324
rect 477862 225200 477984 225328
rect 477548 224880 477644 224992
rect 482160 224896 482216 225008
rect 477552 224274 477648 224396
rect 478646 224236 478702 224358
rect 477552 223786 477648 223892
rect 477862 223776 477984 223904
rect 33176 219357 33382 223223
rect 72954 208656 73584 209538
rect 79331 206980 79685 207942
rect 34939 203662 35194 206806
rect 74345 205038 74614 205722
rect 70812 198094 71316 198850
rect 69048 192402 69552 193032
rect 35539 186862 35794 190006
rect 66150 189252 66780 190008
rect 64545 187664 64831 187864
rect 66801 185801 67014 185968
rect 36139 170062 36394 173206
rect 73332 166446 74088 167202
rect 79506 164178 79884 165312
rect 80892 161532 81522 162036
rect 36739 153262 36994 156406
rect 51408 152838 52794 153468
rect 321100 149336 321500 149736
rect 321183 148391 321445 148653
rect 52164 148226 52220 148371
rect 52724 148226 52780 148370
rect 53284 148226 53340 148370
rect 53844 148217 53900 148370
rect 52500 146702 52556 146848
rect 53060 146702 53116 146848
rect 53620 146702 53676 146848
rect 54180 146702 54236 146848
rect 61334 144890 61390 144966
rect 61684 144816 61740 145040
rect 61908 144900 61964 144956
rect 62356 144816 62412 145040
rect 62580 144900 62636 144956
rect 63028 144816 63084 145040
rect 63252 144900 63308 144956
rect 63700 144816 63756 145040
rect 63924 144900 63980 144956
rect 64372 144816 64428 145040
rect 64596 144900 64652 144956
rect 65044 144816 65100 145040
rect 65268 144900 65324 144956
rect 65716 144816 65772 145040
rect 65940 144900 65996 144956
rect 66388 144816 66444 145040
rect 66612 144900 66668 144956
rect 67060 144816 67116 145040
rect 67284 144900 67340 144956
rect 67732 144816 67788 145040
rect 67956 144900 68012 144956
rect 68404 144816 68460 145040
rect 68628 144900 68684 144956
rect 69076 144816 69132 145040
rect 69300 144900 69356 144956
rect 69748 144816 69804 145040
rect 69972 144900 70028 144956
rect 70420 144816 70476 145040
rect 70644 144900 70700 144956
rect 71092 144816 71148 145040
rect 71316 144900 71372 144956
rect 71764 144816 71820 145040
rect 71988 144900 72044 144956
rect 72436 144816 72492 145040
rect 72660 144900 72716 144956
rect 73108 144816 73164 145040
rect 73332 144900 73388 144956
rect 73780 144816 73836 145040
rect 74004 144900 74060 144956
rect 74452 144816 74508 145040
rect 74676 144900 74732 144956
rect 75124 144816 75180 145040
rect 75348 144900 75404 144956
rect 75796 144816 75852 145040
rect 76020 144900 76076 144956
rect 76468 144816 76524 145040
rect 76692 144900 76748 144956
rect 77140 144816 77196 145040
rect 77364 144900 77420 144956
rect 77812 144816 77868 145040
rect 78036 144900 78092 144956
rect 78484 144816 78540 145040
rect 78708 144900 78764 144956
rect 79156 144816 79212 145040
rect 79380 144900 79436 144956
rect 79828 144816 79884 145040
rect 81270 142380 81648 146412
rect 84422 145174 84478 145361
rect 84663 145226 84797 145302
rect 84870 145174 84926 145361
rect 85111 145226 85245 145302
rect 85318 145174 85374 145361
rect 85559 145226 85693 145302
rect 85990 145166 86046 145353
rect 86231 145226 86365 145302
rect 86662 145166 86718 145353
rect 82494 144633 83152 144978
rect 481908 144704 481964 144816
rect 481908 144144 481964 144256
rect 89264 138432 90720 139328
rect 480410 139324 480466 139446
rect 481908 138096 481964 138208
rect 60984 133560 61362 135828
rect 61908 135380 61964 135436
rect 62244 135268 62300 135546
rect 62580 135380 62636 135436
rect 62916 135268 62972 135546
rect 63252 135380 63308 135436
rect 63588 135268 63644 135546
rect 63924 135380 63980 135436
rect 64260 135268 64316 135546
rect 64596 135380 64652 135436
rect 64932 135268 64988 135546
rect 65268 135380 65324 135436
rect 65604 135268 65660 135546
rect 65940 135380 65996 135436
rect 66276 135268 66332 135546
rect 66612 135380 66668 135436
rect 66948 135268 67004 135546
rect 67284 135380 67340 135436
rect 67620 135268 67676 135546
rect 67956 135380 68012 135436
rect 68292 135268 68348 135546
rect 68628 135268 68684 135546
rect 68964 135380 69020 135436
rect 69188 135380 69244 135436
rect 69636 135268 69692 135546
rect 69860 135380 69916 135436
rect 70308 135268 70364 135546
rect 70532 135380 70588 135436
rect 70980 135268 71036 135546
rect 71204 135380 71260 135436
rect 71652 135268 71708 135546
rect 71876 135380 71932 135436
rect 72324 135268 72380 135546
rect 72548 135380 72604 135436
rect 72996 135268 73052 135546
rect 73220 135380 73276 135436
rect 73668 135268 73724 135546
rect 73892 135380 73948 135436
rect 74340 135268 74396 135546
rect 74564 135380 74620 135436
rect 75012 135268 75068 135546
rect 75236 135380 75292 135436
rect 75684 135268 75740 135546
rect 75908 135380 75964 135436
rect 76356 135268 76412 135546
rect 76580 135380 76636 135436
rect 77028 135268 77084 135546
rect 77252 135380 77308 135436
rect 77700 135268 77756 135546
rect 77924 135380 77980 135436
rect 78372 135268 78428 135546
rect 78596 135380 78652 135436
rect 79044 135268 79100 135546
rect 79268 135380 79324 135436
rect 79716 135268 79772 135546
rect 81270 134946 81648 136458
rect 481376 134952 481472 135058
rect 481690 134934 481812 135062
rect 479906 134444 479962 134566
rect 481376 134444 481472 134566
rect 480158 133956 480214 134078
rect 481380 133956 481476 134078
rect 62132 133262 62188 133411
rect 62692 133262 62748 133411
rect 63252 133262 63308 133411
rect 63812 133262 63868 133411
rect 64372 133257 64428 133416
rect 64932 133257 64988 133416
rect 65492 133257 65548 133416
rect 66052 133257 66108 133416
rect 66612 133257 66668 133416
rect 67172 133257 67228 133416
rect 67732 133257 67788 133416
rect 68292 133257 68348 133416
rect 68852 133257 68908 133416
rect 69412 133257 69468 133416
rect 69972 133257 70028 133416
rect 70532 133257 70588 133416
rect 275900 133100 276500 133700
rect 481380 133520 481476 133626
rect 481690 133510 481812 133638
rect 72314 132174 73070 132804
rect 276069 131825 276331 132087
rect 62748 131040 65646 131292
rect 58556 130697 58620 130947
rect 59960 130683 60016 130853
rect 60353 130736 60409 130906
rect 61755 130683 61811 130853
rect 59780 130447 60083 130503
rect 61577 130445 61880 130502
rect 62748 130158 65646 130410
rect 481908 127904 481964 128016
rect 59850 127386 60102 127638
rect 481908 127344 481964 127456
rect 59115 127082 59193 127246
rect 61110 126630 61866 127008
rect 117460 126788 117516 126844
rect 117684 125780 117740 125836
rect 479150 122488 479206 122610
rect 481908 121296 481964 121408
rect 117908 119844 117964 119900
rect 118132 118948 118188 119004
rect 481376 118152 481472 118258
rect 481690 118134 481812 118262
rect 118356 117940 118412 117996
rect 479654 117730 479710 117852
rect 481376 117730 481472 117852
rect 479402 117120 479458 117242
rect 481380 117120 481476 117242
rect 118580 116932 118636 116988
rect 481380 116720 481476 116826
rect 481690 116710 481812 116838
rect 118804 115924 118860 115980
rect 63513 111275 63569 111371
rect 63875 111368 63931 111474
rect 64889 111196 64945 111352
rect 65143 111308 65199 111556
rect 66033 111275 66089 111371
rect 66395 111368 66451 111474
rect 67409 111196 67465 111352
rect 67663 111308 67719 111556
rect 68553 111275 68609 111371
rect 68915 111368 68971 111474
rect 69929 111196 69985 111352
rect 70183 111308 70239 111556
rect 37674 108612 38556 109620
rect 66906 108738 67536 109116
rect 61468 108515 61636 108571
rect 63850 108503 64165 108559
rect 68152 108469 68212 108581
rect 71008 108500 71450 108556
rect 59598 106974 60606 107352
rect 65898 107226 66528 107604
rect 86412 108538 86640 108738
rect 91476 108738 91728 109620
rect 74340 107352 75096 107856
rect 90468 107478 90846 107856
rect 74074 107016 74196 107072
rect 92484 107352 92988 107856
rect 35188 95508 35244 95584
rect 35524 78102 35580 78178
rect 119028 114916 119084 114972
rect 116564 114020 116620 114076
rect 116340 113012 116396 113068
rect 117236 112004 117292 112060
rect 117460 111444 117516 111500
rect 117684 109988 117740 110044
rect 117908 108448 117964 108504
rect 118132 106992 118188 107048
rect 477383 79083 477645 79345
rect 477300 78000 477700 78400
rect 119264 72760 119904 72820
rect 119264 72600 119904 72660
rect 113274 71442 113904 72072
rect 114660 71694 115164 72198
rect 116067 71564 116239 71620
rect 117470 71614 117534 71802
rect 136072 71442 140860 72828
rect 205006 59033 206669 59840
rect 268506 59472 283122 61362
rect 472600 61200 477800 75600
rect 34600 43200 36200 57600
rect 199200 51600 204464 53800
rect 205440 51600 210800 53800
rect 59800 41100 60400 41700
rect 59983 40083 60245 40345
rect 231800 37200 246200 42200
rect 34992 34128 35048 34184
rect 34362 33876 34418 33932
rect 102400 33800 116800 35400
rect 73422 33624 73478 33680
rect 56538 33372 56594 33428
rect 55404 32624 55460 32680
rect 72162 32624 72218 32680
rect 90180 33120 90236 33176
rect 88920 32624 88976 32680
rect 285400 53400 299800 58600
rect 318083 51883 318345 52145
rect 317900 50500 318500 51100
rect 481418 48922 481474 49044
rect 481908 47712 481964 47824
rect 480683 44683 480945 44945
rect 480500 43100 481100 43700
rect 328104 37548 328230 37604
rect 311346 36328 311472 36384
rect 310886 33078 311014 33200
rect 310896 32768 311002 32864
rect 311346 32768 311472 32864
rect 311976 36084 312102 36140
rect 312310 33078 312438 33200
rect 327686 33078 327814 33200
rect 311976 32764 312102 32860
rect 312328 32764 312434 32860
rect 327696 32768 327802 32864
rect 420714 37304 420840 37360
rect 403956 37060 404082 37116
rect 387072 36816 387198 36872
rect 370314 36572 370440 36628
rect 328104 32768 328230 32864
rect 328734 35840 328860 35896
rect 365526 35596 365652 35652
rect 364896 34630 365022 34686
rect 329110 33078 329238 33200
rect 364486 33078 364614 33200
rect 328734 32764 328860 32860
rect 329128 32764 329234 32860
rect 364496 32768 364602 32864
rect 364896 32768 365022 32864
rect 369040 33348 369152 33404
rect 365910 33078 366038 33200
rect 365526 32764 365652 32860
rect 365928 32764 366034 32860
rect 382284 35352 382410 35408
rect 381654 34378 381780 34434
rect 381286 33078 381414 33200
rect 381296 32768 381402 32864
rect 381654 32768 381780 32864
rect 385840 33348 385952 33404
rect 382710 33078 382838 33200
rect 382284 32764 382410 32860
rect 382728 32764 382834 32860
rect 399168 35108 399294 35164
rect 398538 34126 398664 34182
rect 398086 33078 398214 33200
rect 398096 32768 398202 32864
rect 398538 32768 398664 32864
rect 402640 33348 402752 33404
rect 399510 33078 399638 33200
rect 399168 32764 399294 32860
rect 399528 32764 399634 32860
rect 415926 34924 416052 34980
rect 415296 33874 415422 33930
rect 414886 33078 415014 33200
rect 414896 32768 415002 32864
rect 415296 32768 415422 32864
rect 419440 33348 419552 33404
rect 416310 33078 416438 33200
rect 415926 32764 416052 32860
rect 416328 32764 416434 32860
rect 432820 33078 433812 33200
rect 471492 33606 471618 33662
rect 470288 33348 470400 33404
<< metal2 >>
rect 32228 381332 44128 381388
rect 44240 381332 60928 381388
rect 61040 381332 77728 381388
rect 77840 381332 94528 381388
rect 94640 381332 111328 381388
rect 111440 381332 128128 381388
rect 128240 381332 144928 381388
rect 145040 381332 201712 381388
rect 201824 381332 218512 381388
rect 218624 381332 245280 381388
rect 245392 381332 262080 381388
rect 262192 381332 278880 381388
rect 278992 381332 279104 381388
rect 32228 333424 32284 381332
rect 48344 381220 48384 381276
rect 48496 381220 78708 381276
rect 78764 381220 78804 381276
rect 38152 381108 38192 381164
rect 38304 381108 80052 381164
rect 80108 381108 80148 381164
rect 37480 380996 37520 381052
rect 37632 380996 82628 381052
rect 82684 380996 82724 381052
rect 87460 380994 87470 381086
rect 87560 380994 87920 381086
rect 88032 380994 88068 381086
rect 88564 380968 88592 381060
rect 88704 380968 89066 381060
rect 89156 380968 89170 381060
rect 97644 380994 97662 381086
rect 97752 380994 98112 381086
rect 98224 380994 98260 381086
rect 98756 380968 98784 381060
rect 98896 380968 99258 381060
rect 99348 380968 99372 381060
rect 104260 380994 104270 381086
rect 104360 380994 104720 381086
rect 104832 380994 104868 381086
rect 105364 380968 105392 381060
rect 105504 380968 105866 381060
rect 105956 380968 105970 381060
rect 114444 380994 114462 381086
rect 114552 380994 114912 381086
rect 115024 380994 115060 381086
rect 115556 380968 115584 381060
rect 115696 380968 116058 381060
rect 116148 380968 116172 381060
rect 121060 380994 121070 381086
rect 121160 380994 121520 381086
rect 121632 380994 121668 381086
rect 122164 380968 122192 381060
rect 122304 380968 122666 381060
rect 122756 380968 122770 381060
rect 131244 380994 131262 381086
rect 131352 380994 131712 381086
rect 131824 380994 131860 381086
rect 132356 380968 132384 381060
rect 132496 380968 132858 381060
rect 132948 380968 132972 381060
rect 137860 380994 137870 381086
rect 137960 380994 138320 381086
rect 138432 380994 138468 381086
rect 138964 380968 138992 381060
rect 139104 380968 139466 381060
rect 139556 380968 139570 381060
rect 148044 380994 148062 381086
rect 148152 380994 148512 381086
rect 148624 380994 148660 381086
rect 149156 380968 149184 381060
rect 149296 380968 149658 381060
rect 149748 380968 149772 381060
rect 194660 380994 194670 381086
rect 194760 380994 195120 381086
rect 195232 380994 195268 381086
rect 195764 380968 195792 381060
rect 195904 380968 196266 381060
rect 196356 380968 196370 381060
rect 204844 380994 204862 381086
rect 204952 380994 205312 381086
rect 205424 380994 205460 381086
rect 205956 380968 205984 381060
rect 206096 380968 206458 381060
rect 206548 380968 206572 381060
rect 211460 380994 211470 381086
rect 211560 380994 211920 381086
rect 212032 380994 212068 381086
rect 212564 380968 212592 381060
rect 212704 380968 213066 381060
rect 213156 380968 213170 381060
rect 221644 380994 221662 381086
rect 221752 380994 222112 381086
rect 222224 380994 222260 381086
rect 222756 380968 222784 381060
rect 222896 380968 223258 381060
rect 223348 380968 223372 381060
rect 238260 380994 238270 381086
rect 238360 380994 238720 381086
rect 238832 380994 238868 381086
rect 239364 380968 239392 381060
rect 239504 380968 239866 381060
rect 239956 380968 239970 381060
rect 248444 380994 248462 381086
rect 248552 380994 248912 381086
rect 249024 380994 249060 381086
rect 249556 380968 249584 381060
rect 249696 380968 250058 381060
rect 250148 380968 250172 381060
rect 255060 380994 255070 381086
rect 255160 380994 255520 381086
rect 255632 380994 255668 381086
rect 256164 380968 256192 381060
rect 256304 380968 256666 381060
rect 256756 380968 256770 381060
rect 265244 380994 265262 381086
rect 265352 380994 265712 381086
rect 265824 380994 265860 381086
rect 266356 380968 266384 381060
rect 266496 380968 266858 381060
rect 266948 380968 266972 381060
rect 271860 380994 271870 381086
rect 271960 380994 272320 381086
rect 272432 380994 272468 381086
rect 272964 380968 272992 381060
rect 273104 380968 273466 381060
rect 273556 380968 273570 381060
rect 282044 380994 282062 381086
rect 282152 380994 282512 381086
rect 282624 380994 282660 381086
rect 283156 380968 283184 381060
rect 283296 380968 283658 381060
rect 283748 380968 283772 381060
rect 47672 380884 47712 380940
rect 47824 380884 82740 380940
rect 82796 380884 82836 380940
rect 42968 380772 43008 380828
rect 43120 380772 85428 380828
rect 85484 380772 85524 380828
rect 332100 380778 332806 380830
rect 65144 380660 65184 380716
rect 65296 380660 78820 380716
rect 78876 380660 78916 380716
rect 54952 380548 54992 380604
rect 55104 380548 80164 380604
rect 80220 380548 80260 380604
rect 332100 380602 332154 380778
rect 33462 380400 34702 380490
rect 54280 380436 54320 380492
rect 54432 380436 82516 380492
rect 82572 380436 82612 380492
rect 87394 380458 87450 380602
rect 87582 380458 89040 380602
rect 89172 380458 97642 380602
rect 97774 380458 99232 380602
rect 99364 380458 104250 380602
rect 104382 380458 105840 380602
rect 105972 380458 114442 380602
rect 114574 380458 116032 380602
rect 116164 380458 121050 380602
rect 121182 380458 122640 380602
rect 122772 380458 131242 380602
rect 131374 380458 132832 380602
rect 132964 380458 137850 380602
rect 137982 380458 139440 380602
rect 139572 380458 148042 380602
rect 148174 380458 149632 380602
rect 149764 380458 194650 380602
rect 194782 380458 196240 380602
rect 196372 380458 204842 380602
rect 204974 380458 206432 380602
rect 206564 380458 211450 380602
rect 211582 380458 213040 380602
rect 213172 380458 221642 380602
rect 221774 380458 223232 380602
rect 223364 380458 238250 380602
rect 238382 380458 239840 380602
rect 239972 380458 248442 380602
rect 248574 380458 250032 380602
rect 250164 380458 255050 380602
rect 255182 380458 256640 380602
rect 256772 380458 265242 380602
rect 265374 380458 266832 380602
rect 266964 380458 271850 380602
rect 271982 380458 273440 380602
rect 273572 380458 282042 380602
rect 282174 380458 283632 380602
rect 283764 380458 332154 380602
rect 33462 366000 33600 380400
rect 34600 366000 34702 380400
rect 64472 380324 64512 380380
rect 64624 380324 82852 380380
rect 82908 380324 82948 380380
rect 59768 380212 59808 380268
rect 59920 380212 85652 380268
rect 85708 380212 85748 380268
rect 332100 380250 332154 380458
rect 332744 380250 332806 380778
rect 332100 380188 332806 380250
rect 77078 380100 77110 380156
rect 77228 380100 78932 380156
rect 78988 380100 81984 380156
rect 82096 380100 82110 380156
rect 71752 379988 71792 380044
rect 71904 379988 80276 380044
rect 80332 379988 80372 380044
rect 71080 379876 71120 379932
rect 71232 379876 82404 379932
rect 82460 379876 82500 379932
rect 77754 379764 77784 379820
rect 77898 379764 81312 379820
rect 81424 379764 82964 379820
rect 83020 379764 83060 379820
rect 76568 379652 76608 379708
rect 76720 379652 85876 379708
rect 85932 379652 85964 379708
rect 79004 379540 79044 379596
rect 79100 379540 98784 379596
rect 98896 379540 98936 379596
rect 80348 379428 80388 379484
rect 80444 379428 88592 379484
rect 88704 379428 88744 379484
rect 82252 379316 82292 379372
rect 82348 379316 87920 379372
rect 88032 379316 88072 379372
rect 83036 379204 83076 379260
rect 83132 379204 98112 379260
rect 98224 379204 98264 379260
rect 79116 379092 79156 379148
rect 79212 379092 115584 379148
rect 115696 379092 115736 379148
rect 80460 378980 80500 379036
rect 80556 378980 105392 379036
rect 105504 378980 105520 379036
rect 82140 378868 82180 378924
rect 82236 378868 104720 378924
rect 104832 378868 104857 378924
rect 83148 378756 83188 378812
rect 83244 378756 114912 378812
rect 115024 378756 115064 378812
rect 37060 378594 37070 378686
rect 37160 378594 37520 378686
rect 37632 378594 37668 378686
rect 38164 378568 38192 378660
rect 38304 378568 38666 378660
rect 38756 378568 38770 378660
rect 47244 378594 47262 378686
rect 47352 378594 47712 378686
rect 47824 378594 47860 378686
rect 48356 378568 48384 378660
rect 48496 378568 48858 378660
rect 48948 378568 48972 378660
rect 53860 378594 53870 378686
rect 53960 378594 54320 378686
rect 54432 378594 54468 378686
rect 54964 378568 54992 378660
rect 55104 378568 55466 378660
rect 55556 378568 55570 378660
rect 64044 378594 64062 378686
rect 64152 378594 64512 378686
rect 64624 378594 64660 378686
rect 65156 378568 65184 378660
rect 65296 378568 65658 378660
rect 65748 378568 65772 378660
rect 70660 378594 70670 378686
rect 70760 378594 71120 378686
rect 71232 378594 71268 378686
rect 71764 378568 71792 378660
rect 71904 378568 72266 378660
rect 72356 378568 72370 378660
rect 76644 378594 76662 378686
rect 76752 378594 77112 378686
rect 77224 378594 77260 378686
rect 77756 378568 77784 378660
rect 77896 378568 78258 378660
rect 78348 378568 78372 378660
rect 79228 378644 79268 378700
rect 79324 378644 132384 378700
rect 132496 378644 132536 378700
rect 80572 378532 80612 378588
rect 80668 378532 122192 378588
rect 122304 378532 122344 378588
rect 82028 378420 82068 378476
rect 82124 378420 121520 378476
rect 121632 378420 121672 378476
rect 83260 378308 83300 378364
rect 83356 378308 131712 378364
rect 131824 378308 131864 378364
rect 35518 378058 35550 378202
rect 35872 378058 37050 378202
rect 37182 378058 38640 378202
rect 38772 378058 47242 378202
rect 47374 378058 48832 378202
rect 48964 378058 53850 378202
rect 53982 378058 55440 378202
rect 55572 378058 64042 378202
rect 64174 378058 65632 378202
rect 65764 378058 70650 378202
rect 70782 378058 72240 378202
rect 72372 378058 76642 378202
rect 76774 378058 78232 378202
rect 78364 378058 78438 378202
rect 79340 378196 79380 378252
rect 79436 378196 149184 378252
rect 149296 378196 149336 378252
rect 80684 378084 80724 378140
rect 80780 378084 138992 378140
rect 139104 378084 139144 378140
rect 81916 377972 81956 378028
rect 82012 377972 138320 378028
rect 138432 377972 138472 378028
rect 83372 377860 83412 377916
rect 83468 377860 148512 377916
rect 148624 377860 148664 377916
rect 79452 377748 79492 377804
rect 79548 377748 205984 377804
rect 206096 377748 206136 377804
rect 80796 377636 80836 377692
rect 80892 377636 195792 377692
rect 195904 377636 195944 377692
rect 81804 377524 81844 377580
rect 81900 377524 195120 377580
rect 195232 377524 195272 377580
rect 83484 377412 83524 377468
rect 83580 377412 205312 377468
rect 205424 377412 205464 377468
rect 79564 377300 79604 377356
rect 79660 377300 222784 377356
rect 222896 377300 222936 377356
rect 80908 377188 80948 377244
rect 81004 377188 212592 377244
rect 212704 377188 212744 377244
rect 81692 377076 81732 377132
rect 81788 377076 211920 377132
rect 212032 377076 212072 377132
rect 83596 376964 83636 377020
rect 83692 376964 222112 377020
rect 222224 376964 222264 377020
rect 79676 376852 79716 376908
rect 79772 376852 249584 376908
rect 249696 376852 249736 376908
rect 81020 376740 81060 376796
rect 81116 376740 239392 376796
rect 239504 376740 239544 376796
rect 81580 376628 81620 376684
rect 81676 376628 238720 376684
rect 238832 376628 238872 376684
rect 83708 376516 83748 376572
rect 83804 376516 248912 376572
rect 249024 376516 249064 376572
rect 79788 376404 79828 376460
rect 79884 376404 266384 376460
rect 266496 376404 266536 376460
rect 81132 376292 81172 376348
rect 81228 376292 256192 376348
rect 256304 376292 256344 376348
rect 81468 376180 81508 376236
rect 81564 376180 255520 376236
rect 255632 376180 255672 376236
rect 83820 376068 83860 376124
rect 83916 376068 265712 376124
rect 265824 376068 265864 376124
rect 79900 375956 79940 376012
rect 79996 375956 283184 376012
rect 283296 375956 283336 376012
rect 81244 375844 81284 375900
rect 81340 375844 272992 375900
rect 273104 375844 273144 375900
rect 427200 375800 442000 376000
rect 81356 375732 81396 375788
rect 81452 375732 272320 375788
rect 272432 375732 272472 375788
rect 83932 375620 83972 375676
rect 84028 375620 282512 375676
rect 282624 375620 282664 375676
rect 93380 374927 93436 374976
rect 78708 373072 78764 373184
rect 68964 370786 69020 370826
rect 68852 370542 68908 370582
rect 63378 367542 64890 367668
rect 63378 366912 63504 367542
rect 64764 366912 64890 367542
rect 63378 366786 64890 366912
rect 33462 365904 34702 366000
rect 68292 366150 68348 366190
rect 33492 363600 34716 363688
rect 33492 349200 33600 363600
rect 34600 349200 34716 363600
rect 68068 362246 68124 362286
rect 66024 361620 66906 361746
rect 65268 360864 65772 360990
rect 65268 360360 65394 360864
rect 65646 360360 65772 360864
rect 65268 360234 65772 360360
rect 66024 360360 66150 361620
rect 66780 360360 66906 361620
rect 66024 360234 66906 360360
rect 63478 360122 63542 360149
rect 64762 360116 64778 360172
rect 64940 360116 65106 360172
rect 63478 359215 63542 359934
rect 46705 359151 63542 359215
rect 64092 359549 64148 359581
rect 46705 357270 46765 359151
rect 63000 358470 63504 358596
rect 64092 358554 64148 359493
rect 63000 358092 63126 358470
rect 63378 358092 63504 358470
rect 63632 358418 63662 358494
rect 63798 358418 63822 358494
rect 63000 357966 63504 358092
rect 63693 357782 63769 358418
rect 64764 359325 64820 359365
rect 64764 358554 64820 359269
rect 65050 359101 65106 360116
rect 68068 359549 68124 362190
rect 68068 359453 68124 359493
rect 68292 359325 68348 366094
rect 68292 359229 68348 359269
rect 68516 365662 68572 365702
rect 65050 359020 65106 359045
rect 68516 359101 68572 365606
rect 68516 359005 68572 359045
rect 68740 364442 68796 364482
rect 64304 358418 64332 358494
rect 64472 358418 64496 358494
rect 64092 358341 64148 358367
rect 49277 357706 63769 357782
rect 49277 357270 49337 357706
rect 64365 357644 64441 358418
rect 64764 358350 64820 358367
rect 64365 357588 68572 357644
rect 64365 357242 64441 357588
rect 33492 349086 34716 349200
rect 32808 338132 32900 338156
rect 32808 337680 32900 338042
rect 32808 337540 32900 337568
rect 33226 338148 33370 338222
rect 32782 337120 32874 337156
rect 32782 336648 32874 337008
rect 32782 336540 32874 336558
rect 33226 336670 33370 338016
rect 33226 336260 33370 336538
rect 34020 337680 34076 337720
rect 33078 336226 33506 336260
rect 33078 335888 33120 336226
rect 33462 335888 33506 336226
rect 33078 335846 33506 335888
rect 32228 316624 32284 333312
rect 32808 327940 32900 327964
rect 32808 327488 32900 327850
rect 32808 327348 32900 327376
rect 33226 327956 33370 335846
rect 32782 326816 32874 326852
rect 32782 326344 32874 326704
rect 32782 326236 32874 326254
rect 33226 326366 33370 327824
rect 32808 321332 32900 321356
rect 32808 320880 32900 321242
rect 32808 320740 32900 320768
rect 33226 321348 33370 326234
rect 32782 320320 32874 320356
rect 32782 319848 32874 320208
rect 32782 319740 32874 319758
rect 33226 319870 33370 321216
rect 32228 299824 32284 316512
rect 32808 311140 32900 311164
rect 32808 310688 32900 311050
rect 32808 310548 32900 310576
rect 33226 311156 33370 319738
rect 32782 310016 32874 310052
rect 32782 309544 32874 309904
rect 32782 309436 32874 309454
rect 33226 309566 33370 311024
rect 33226 309060 33370 309434
rect 32108 288326 32164 288368
rect 32108 287280 32164 288270
rect 32108 287136 32164 287168
rect 32228 283024 32284 299712
rect 32358 308964 33370 309060
rect 33460 320880 33516 320920
rect 32358 304556 32454 308964
rect 32430 304430 32454 304556
rect 32358 302962 32454 304430
rect 32566 304526 32632 304563
rect 32566 304080 32632 304462
rect 32566 303942 32632 303968
rect 32900 304080 32956 304120
rect 32438 302836 32454 302962
rect 32358 294244 32454 302836
rect 32540 303520 32612 303544
rect 32540 302936 32612 303408
rect 32540 302826 32612 302860
rect 32448 294118 32454 294244
rect 32358 292650 32454 294118
rect 32562 294224 32630 294240
rect 32562 293888 32630 294140
rect 32562 293744 32630 293776
rect 32434 292524 32454 292650
rect 32540 293216 32610 293240
rect 32540 292630 32610 293104
rect 32540 292534 32610 292546
rect 32358 288694 32454 292524
rect 32358 287904 32454 288570
rect 32570 288670 32656 288682
rect 32570 288326 32656 288596
rect 32570 288246 32656 288270
rect 32446 287776 32454 287904
rect 32358 287574 32454 287776
rect 32554 287882 32628 287896
rect 32340 287280 32396 287337
rect 32340 284284 32396 287168
rect 32554 286768 32628 287804
rect 32554 286720 32732 286768
rect 32628 286608 32676 286720
rect 32554 286586 32732 286608
rect 32676 285628 32732 286586
rect 32676 285532 32732 285572
rect 32788 286412 32844 286452
rect 32564 285180 32620 285220
rect 32340 284188 32396 284228
rect 32452 284732 32508 284772
rect 32228 275772 32284 282912
rect 32452 277088 32508 284676
rect 32452 276936 32508 276976
rect 32564 276416 32620 285124
rect 32788 281904 32844 286356
rect 32900 284396 32956 303968
rect 33236 303520 33292 303560
rect 33012 293888 33068 293928
rect 33012 284844 33068 293776
rect 33124 293216 33180 293256
rect 33124 285292 33180 293104
rect 33236 285740 33292 303408
rect 33348 298704 33404 298744
rect 33348 286300 33404 298592
rect 33348 286204 33404 286244
rect 33236 285644 33292 285684
rect 33124 285196 33180 285236
rect 33012 284748 33068 284788
rect 33460 284508 33516 320768
rect 33796 320320 33852 320360
rect 33572 310688 33628 310728
rect 33572 284956 33628 310576
rect 33684 310016 33740 310056
rect 33684 285404 33740 309904
rect 33796 285852 33852 320208
rect 33908 315504 33964 315544
rect 33908 286188 33964 315392
rect 33908 286092 33964 286132
rect 33796 285756 33852 285796
rect 33684 285308 33740 285348
rect 33572 284860 33628 284900
rect 34020 284620 34076 337568
rect 34356 337120 34412 337160
rect 46705 337094 46765 337354
rect 49277 337090 49337 337350
rect 34132 327488 34188 327528
rect 34132 285068 34188 327376
rect 34244 326816 34300 326856
rect 34244 285516 34300 326704
rect 34356 285964 34412 337008
rect 34580 337036 34636 337046
rect 34468 332304 34524 332344
rect 34468 286076 34524 332192
rect 34468 285980 34524 286020
rect 34356 285868 34412 285908
rect 34244 285420 34300 285460
rect 34132 284972 34188 285012
rect 34020 284524 34076 284564
rect 33460 284412 33516 284452
rect 32900 284300 32956 284340
rect 32788 281752 32844 281792
rect 33526 283874 33670 283902
rect 33108 277540 33200 277564
rect 33108 277088 33200 277450
rect 33108 276948 33200 276976
rect 33526 277556 33670 283714
rect 32564 276264 32620 276304
rect 33082 276416 33174 276452
rect 33082 275944 33174 276304
rect 33082 275836 33174 275854
rect 33526 275966 33670 277424
rect 32228 275716 32606 275772
rect 32550 122424 32606 275716
rect 33526 275648 33670 275834
rect 33695 257206 34047 257276
rect 33695 254062 33739 257206
rect 33994 254062 34047 257206
rect 33695 254010 34047 254062
rect 34580 241276 34636 336980
rect 68516 337036 68572 357588
rect 68516 336970 68572 336980
rect 36486 335212 36546 335472
rect 36726 335216 36786 335476
rect 39271 335208 39331 335468
rect 41151 335208 41211 335468
rect 41326 335216 41386 335476
rect 44138 335340 44198 335600
rect 46871 335330 46931 335590
rect 47959 335336 48019 335596
rect 49047 335332 49107 335592
rect 50135 335324 50195 335584
rect 65688 335220 65748 335516
rect 65868 335220 65928 335516
rect 66048 335220 66108 335516
rect 66228 335220 66288 335516
rect 66408 335220 66468 335516
rect 36486 313966 36546 315308
rect 36726 315085 36786 315265
rect 36726 315015 36786 315029
rect 39271 314616 39331 315280
rect 41151 314966 41211 315255
rect 41151 314895 41211 314906
rect 41326 314729 41386 315268
rect 44138 315085 44198 315389
rect 44138 315009 44198 315029
rect 46265 314966 46325 314984
rect 41326 314656 41386 314673
rect 42308 314841 42364 314864
rect 36486 313896 36546 313906
rect 39200 314556 39331 314616
rect 35028 313488 36036 313614
rect 35028 312984 35154 313488
rect 35910 312984 36036 313488
rect 38396 313604 38596 313616
rect 38396 313329 38413 313604
rect 38578 313329 38596 313604
rect 39200 313339 39260 314556
rect 41725 313623 41985 313646
rect 39872 313597 40072 313616
rect 38396 313314 38596 313329
rect 39872 313333 39889 313597
rect 40051 313333 40072 313597
rect 41725 313357 41744 313623
rect 41962 313357 41985 313623
rect 41725 313338 41985 313357
rect 39872 313314 40072 313333
rect 35028 312858 36036 312984
rect 42308 310664 42364 314785
rect 41668 310608 42364 310664
rect 42532 314617 42588 314643
rect 42532 309724 42588 314561
rect 42714 313614 43344 313740
rect 42714 312858 42840 313614
rect 43218 312858 43344 313614
rect 43974 313687 44478 313740
rect 43974 313488 44030 313687
rect 43596 313428 44030 313488
rect 44407 313428 44478 313687
rect 43596 313362 44478 313428
rect 45447 313601 45647 313624
rect 45447 313339 45467 313601
rect 45631 313339 45647 313601
rect 45447 313322 45647 313339
rect 46265 313330 46325 314906
rect 46871 314729 46931 315387
rect 46871 314651 46931 314673
rect 47959 314729 48019 315387
rect 49047 315122 49107 315402
rect 50135 315118 50195 315392
rect 65688 315130 65748 315268
rect 65868 315130 65928 315268
rect 47959 314651 48019 314673
rect 62343 315084 62400 315094
rect 49364 314413 49420 314453
rect 48764 313634 49026 313649
rect 46923 313610 47123 313624
rect 46923 313336 46935 313610
rect 47111 313336 47123 313610
rect 48764 313364 48779 313634
rect 49011 313364 49026 313634
rect 48764 313345 49026 313364
rect 46923 313322 47123 313336
rect 42714 312732 43344 312858
rect 42714 310842 43344 310968
rect 42714 310338 42840 310842
rect 43218 310338 43344 310842
rect 49364 310664 49420 314357
rect 48713 310608 49420 310664
rect 49588 314189 49644 314229
rect 42714 310212 43344 310338
rect 49588 309724 49644 314133
rect 60228 313362 61362 313488
rect 60228 313110 60354 313362
rect 61236 313110 61362 313362
rect 60228 312984 61362 313110
rect 56644 312173 56700 312183
rect 56644 311696 56700 312117
rect 60228 311850 61362 311976
rect 60228 311220 60354 311850
rect 61236 311220 61362 311850
rect 62343 311514 62400 315027
rect 65750 315035 65826 315062
rect 62692 313964 62748 314006
rect 62692 313012 62748 313908
rect 64135 313964 64192 313974
rect 63084 313741 63140 313751
rect 63084 313073 63140 313685
rect 62624 312956 62636 313012
rect 62804 312956 62819 313012
rect 63084 312859 63140 312886
rect 62734 311525 62798 311544
rect 62343 311457 62734 311514
rect 62734 311316 62798 311337
rect 64135 311457 64192 313907
rect 64386 312732 65520 312858
rect 64386 312480 64512 312732
rect 65394 312480 65520 312732
rect 64386 312354 65520 312480
rect 64135 311266 64192 311287
rect 64520 311555 64596 311599
rect 64520 311307 64526 311555
rect 64590 311307 64596 311555
rect 60228 311094 61362 311220
rect 64184 311165 64240 311184
rect 49896 310842 50526 310968
rect 49896 310338 50022 310842
rect 50400 310338 50526 310842
rect 64184 310842 64240 311041
rect 64184 310703 64240 310716
rect 49896 310212 50526 310338
rect 52708 310598 52947 310664
rect 64520 310611 64596 311307
rect 64520 310520 64596 310535
rect 41710 309668 42588 309724
rect 48748 309668 49644 309724
rect 50526 309582 51408 309708
rect 50526 309078 50652 309582
rect 51282 309078 51408 309582
rect 50526 308952 51408 309078
rect 52708 308767 52947 310398
rect 57886 310424 58126 310447
rect 57886 310206 57903 310424
rect 58105 310206 58126 310424
rect 57886 310183 58126 310206
rect 58464 309582 58968 309708
rect 58464 308952 58590 309582
rect 58842 308952 58968 309582
rect 58464 308826 58968 308952
rect 52708 308464 52947 308528
rect 53871 308460 53900 308560
rect 54100 308460 65584 308560
rect 51610 308285 62680 308297
rect 51610 308134 51619 308285
rect 51968 308134 62680 308285
rect 51610 308124 62680 308134
rect 51636 307696 51956 308124
rect 62604 307669 62680 308124
rect 65508 307776 65584 308460
rect 65750 307728 65826 314979
rect 66048 315035 66108 315260
rect 66048 314961 66108 314979
rect 66228 315035 66288 315273
rect 66228 314961 66288 314979
rect 65927 313517 65984 313542
rect 65927 311457 65984 313461
rect 66408 312017 66468 315308
rect 66320 311957 66468 312017
rect 67719 313293 67776 313333
rect 66320 311576 66380 311957
rect 66320 311425 66380 311445
rect 67719 311457 67776 313237
rect 68740 312173 68796 364386
rect 68852 314861 68908 370486
rect 68852 314765 68908 314805
rect 68964 314637 69020 370730
rect 68964 314541 69020 314581
rect 69076 369322 69132 369362
rect 69076 314413 69132 369266
rect 69076 314317 69132 314357
rect 69188 369078 69244 369118
rect 69188 314189 69244 369022
rect 69188 314093 69244 314133
rect 69300 365418 69356 365458
rect 69300 313965 69356 365362
rect 69636 364930 69692 364956
rect 69524 364686 69580 364706
rect 69300 313869 69356 313909
rect 69412 362490 69468 362530
rect 69412 313741 69468 362434
rect 69412 313636 69468 313685
rect 69524 313517 69580 364630
rect 69524 313421 69580 313461
rect 69636 313293 69692 364874
rect 74452 364198 74508 364223
rect 71652 363954 71708 363994
rect 71540 363710 71596 363750
rect 71428 363466 71484 363506
rect 71316 361758 71372 361798
rect 69636 313197 69692 313237
rect 69748 357122 69804 357162
rect 68740 312077 68796 312117
rect 65927 311266 65984 311287
rect 67719 311266 67776 311287
rect 68544 311220 69552 311346
rect 65976 311165 66032 311184
rect 65976 310842 66032 311041
rect 65976 310703 66032 310716
rect 67768 311165 67824 311184
rect 67768 310842 67824 311041
rect 68544 310968 68670 311220
rect 69426 310968 69552 311220
rect 68544 310842 69552 310968
rect 67768 310703 67824 310716
rect 67446 310611 67522 310640
rect 67446 307760 67522 310535
rect 68976 310414 69088 310464
rect 68976 284032 69088 310214
rect 37707 282078 38635 282086
rect 37707 281653 37740 282078
rect 38303 281653 38635 282078
rect 37707 281651 38635 281653
rect 37535 249473 38644 249485
rect 37535 248893 37590 249473
rect 38138 248893 38644 249473
rect 37535 248888 38644 248893
rect 58464 247968 59346 248094
rect 58464 247086 58590 247968
rect 59220 247086 59346 247968
rect 58464 245622 59346 247086
rect 56196 245322 59346 245622
rect 60102 246330 60982 246456
rect 60102 245448 60228 246330
rect 60858 245448 60982 246330
rect 60102 245262 60982 245448
rect 56196 244962 60982 245262
rect 63756 244692 64764 244818
rect 63756 243936 63882 244692
rect 64638 243936 64764 244692
rect 63756 243882 64764 243936
rect 46116 243784 46172 243824
rect 34580 241220 35084 241276
rect 34295 240406 34647 240476
rect 34295 237262 34339 240406
rect 34594 237262 34647 240406
rect 34295 237210 34647 237262
rect 33126 223223 33425 223279
rect 33126 219357 33176 223223
rect 33382 219357 33425 223223
rect 33126 219314 33425 219357
rect 35028 207564 35084 241220
rect 46116 240872 46172 243728
rect 64036 243784 64092 243796
rect 46116 240776 46172 240816
rect 47908 243662 47964 243702
rect 47908 240750 47964 243606
rect 62244 243662 62300 243718
rect 47908 240654 47964 240694
rect 49700 243540 49756 243580
rect 49700 240628 49756 243484
rect 60452 243540 60508 243584
rect 49700 240532 49756 240572
rect 51492 243418 51548 243458
rect 51492 240506 51548 243362
rect 58660 243418 58716 243450
rect 51492 240410 51548 240450
rect 53284 243296 53340 243336
rect 53284 240384 53340 243240
rect 56868 243296 56924 243338
rect 53284 240288 53340 240328
rect 55076 243174 55132 243196
rect 55076 240262 55132 243118
rect 55076 240166 55132 240206
rect 56868 240140 56924 243240
rect 56868 240044 56924 240084
rect 49839 240030 50439 240031
rect 49644 239904 51786 240030
rect 58660 240018 58716 243362
rect 58660 239922 58716 239962
rect 49644 239778 49770 239904
rect 51660 239778 51786 239904
rect 60452 239896 60508 243484
rect 60452 239800 60508 239840
rect 49644 239652 51786 239778
rect 62244 239774 62300 243606
rect 62244 239678 62300 239718
rect 64036 239652 64092 243728
rect 67158 243180 68040 243306
rect 67158 242298 67284 243180
rect 67914 242298 68040 243180
rect 67158 242172 68040 242298
rect 65638 241794 67024 241920
rect 65638 241290 65764 241794
rect 66898 241290 67024 241794
rect 65638 241164 67024 241290
rect 49839 239304 50439 239652
rect 64036 239556 64092 239596
rect 37707 237878 39933 237886
rect 37707 237453 37740 237878
rect 38303 237453 39933 237878
rect 37707 237451 39933 237453
rect 68976 234773 69088 283922
rect 68976 234523 69088 234573
rect 64827 233982 64849 234149
rect 65109 233982 66949 234149
rect 69748 233996 69804 357066
rect 69636 233940 69804 233996
rect 69860 356878 69916 356918
rect 69860 233996 69916 356822
rect 70084 356634 70140 356674
rect 69972 356390 70028 356430
rect 69972 235676 70028 356334
rect 70084 235788 70140 356578
rect 71204 353706 71260 353746
rect 71092 353462 71148 353502
rect 70980 353218 71036 353258
rect 70868 352974 70924 353014
rect 70756 352730 70812 352770
rect 70644 352486 70700 352526
rect 70532 352242 70588 352282
rect 70420 351998 70476 352038
rect 70308 351754 70364 351794
rect 70196 351510 70252 351550
rect 70196 235900 70252 351454
rect 70308 236012 70364 351698
rect 70420 236124 70476 351942
rect 70532 236236 70588 352186
rect 70644 236348 70700 352430
rect 70756 236460 70812 352674
rect 70868 236572 70924 352918
rect 70980 236684 71036 353162
rect 71092 236796 71148 353406
rect 71204 236908 71260 353650
rect 71316 237020 71372 361702
rect 71428 237132 71484 363410
rect 71540 237244 71596 363654
rect 71652 237356 71708 363898
rect 73220 363222 73276 363262
rect 73108 362978 73164 363018
rect 72996 362734 73052 362774
rect 72884 361514 72940 361554
rect 71764 351266 71820 351306
rect 71764 237468 71820 351210
rect 71876 351022 71932 351062
rect 71876 237580 71932 350966
rect 71988 350778 72044 350818
rect 71988 237692 72044 350722
rect 72100 350534 72156 350574
rect 72100 237804 72156 350478
rect 72212 350290 72268 350330
rect 72212 237916 72268 350234
rect 72324 350046 72380 350086
rect 72324 238028 72380 349990
rect 72436 349802 72492 349842
rect 72436 238140 72492 349746
rect 72548 349558 72604 349598
rect 72548 238252 72604 349502
rect 72660 349314 72716 349354
rect 72660 238364 72716 349258
rect 72772 349070 72828 349110
rect 72772 238476 72828 349014
rect 72884 238588 72940 361458
rect 72996 238700 73052 362678
rect 73108 238812 73164 362922
rect 73220 238924 73276 363166
rect 73332 356146 73388 356186
rect 73332 240872 73388 356090
rect 73332 240776 73388 240816
rect 73444 355902 73500 355942
rect 73444 240750 73500 355846
rect 73444 240654 73500 240694
rect 73556 355658 73612 355698
rect 73556 240628 73612 355602
rect 73556 240532 73612 240572
rect 73668 355414 73724 355454
rect 73668 240506 73724 355358
rect 73668 240410 73724 240450
rect 73780 355170 73836 355210
rect 73780 240384 73836 355114
rect 73780 240288 73836 240328
rect 73892 354926 73948 354966
rect 73892 240262 73948 354870
rect 73892 240166 73948 240206
rect 74004 354682 74060 354722
rect 74004 240140 74060 354626
rect 74004 240044 74060 240084
rect 74116 354438 74172 354478
rect 74116 240018 74172 354382
rect 74116 239922 74172 239962
rect 74228 354194 74284 354234
rect 74228 239896 74284 354138
rect 74228 239800 74284 239840
rect 74340 353950 74396 353990
rect 74340 239774 74396 353894
rect 74340 239678 74396 239718
rect 74452 239652 74508 364142
rect 78708 336812 78764 372624
rect 77364 336756 78764 336812
rect 78820 373072 78876 373184
rect 76356 285964 76412 286004
rect 76244 285852 76300 285892
rect 76132 285740 76188 285780
rect 76020 285628 76076 285668
rect 75908 285516 75964 285556
rect 75796 285404 75852 285444
rect 75684 285292 75740 285332
rect 75572 285180 75628 285220
rect 75460 285068 75516 285108
rect 75348 284956 75404 284996
rect 75236 284844 75292 284884
rect 75124 284732 75180 284772
rect 75012 284620 75068 284660
rect 74900 284508 74956 284548
rect 74788 284396 74844 284436
rect 74676 284284 74732 284324
rect 74676 245492 74732 284228
rect 74788 245736 74844 284340
rect 74900 245980 74956 284452
rect 75012 246224 75068 284564
rect 75124 249396 75180 284676
rect 75236 249640 75292 284788
rect 75348 249884 75404 284900
rect 75460 250128 75516 285012
rect 75572 256960 75628 285124
rect 75572 256864 75628 256904
rect 75684 256716 75740 285236
rect 75684 256620 75740 256660
rect 75796 256472 75852 285348
rect 75796 256376 75852 256416
rect 75908 256228 75964 285460
rect 76020 257204 76076 285572
rect 76132 257448 76188 285684
rect 76244 257692 76300 285796
rect 76356 257936 76412 285908
rect 76356 257840 76412 257880
rect 76244 257596 76300 257636
rect 76132 257352 76188 257392
rect 76020 257108 76076 257148
rect 75908 256132 75964 256172
rect 75460 250032 75516 250072
rect 75348 249788 75404 249828
rect 75236 249544 75292 249584
rect 75124 249300 75180 249340
rect 77364 246468 77420 336756
rect 78820 336700 78876 372624
rect 77476 336644 78876 336700
rect 78932 373072 78988 373184
rect 77476 246712 77532 336644
rect 78932 336588 78988 372624
rect 77588 336532 78988 336588
rect 79044 373072 79100 373184
rect 77588 246956 77644 336532
rect 79044 336476 79100 372624
rect 77700 336420 79100 336476
rect 79156 373072 79212 373184
rect 77700 247200 77756 336420
rect 79156 336364 79212 372624
rect 77812 336308 79212 336364
rect 79268 373072 79324 373184
rect 77812 247444 77868 336308
rect 79268 336252 79324 372624
rect 77924 336196 79324 336252
rect 79380 373072 79436 373184
rect 77924 247688 77980 336196
rect 79380 336140 79436 372624
rect 78036 336084 79436 336140
rect 79492 373072 79548 373184
rect 78036 247932 78092 336084
rect 79492 336028 79548 372624
rect 78148 335972 79548 336028
rect 79604 373072 79660 373184
rect 78148 248176 78204 335972
rect 79604 335916 79660 372624
rect 78260 335860 79660 335916
rect 79716 373072 79772 373184
rect 78260 248420 78316 335860
rect 79716 335804 79772 372624
rect 78372 335748 79772 335804
rect 79828 373072 79884 373184
rect 78372 248664 78428 335748
rect 79828 335692 79884 372624
rect 78484 335636 79884 335692
rect 79940 373072 79996 373184
rect 78484 248908 78540 335636
rect 79940 335580 79996 372624
rect 78596 335524 79996 335580
rect 80052 373072 80108 373184
rect 78596 249152 78652 335524
rect 80052 335468 80108 372624
rect 78708 335412 80108 335468
rect 80164 373072 80220 373184
rect 78708 250372 78764 335412
rect 80164 335356 80220 372624
rect 78820 335300 80220 335356
rect 80276 373072 80332 373184
rect 78820 250616 78876 335300
rect 80276 335244 80332 372624
rect 78932 335188 80332 335244
rect 80388 373072 80444 373184
rect 78932 250860 78988 335188
rect 80388 335132 80444 372624
rect 79044 335076 80444 335132
rect 80500 373072 80556 373184
rect 79044 251104 79100 335076
rect 80500 335020 80556 372624
rect 79156 334964 80556 335020
rect 80612 373072 80668 373184
rect 79156 251348 79212 334964
rect 80612 334908 80668 372624
rect 79268 334852 80668 334908
rect 80724 373072 80780 373184
rect 79268 251592 79324 334852
rect 80724 334796 80780 372624
rect 79380 334740 80780 334796
rect 80836 373072 80892 373184
rect 79380 251836 79436 334740
rect 80836 334684 80892 372624
rect 79492 334628 80892 334684
rect 80948 373072 81004 373184
rect 79492 252080 79548 334628
rect 80948 334572 81004 372624
rect 79604 334516 81004 334572
rect 81060 373072 81116 373184
rect 79604 252324 79660 334516
rect 81060 334460 81116 372624
rect 79716 334404 81116 334460
rect 81172 373072 81228 373184
rect 79716 252568 79772 334404
rect 81172 334348 81228 372624
rect 79828 334292 81228 334348
rect 81284 373072 81340 373184
rect 79828 252812 79884 334292
rect 81284 334236 81340 372624
rect 79940 334180 81340 334236
rect 81396 373072 81452 373184
rect 79940 253056 79996 334180
rect 81396 334124 81452 372624
rect 80052 334068 81452 334124
rect 81508 373072 81564 373184
rect 80052 253300 80108 334068
rect 81508 334012 81564 372624
rect 80164 333956 81564 334012
rect 81620 373072 81676 373184
rect 80164 253544 80220 333956
rect 81620 333900 81676 372624
rect 80276 333844 81676 333900
rect 81732 373072 81788 373184
rect 80276 253788 80332 333844
rect 81732 333788 81788 372624
rect 80388 333732 81788 333788
rect 81844 373072 81900 373184
rect 80388 254032 80444 333732
rect 81844 333676 81900 372624
rect 80500 333620 81900 333676
rect 81956 373072 82012 373184
rect 80500 254276 80556 333620
rect 81956 333564 82012 372624
rect 80612 333508 82012 333564
rect 82068 373072 82124 373184
rect 80612 254520 80668 333508
rect 82068 333452 82124 372624
rect 80724 333396 82124 333452
rect 82180 373072 82236 373184
rect 80724 254764 80780 333396
rect 82180 333340 82236 372624
rect 80836 333284 82236 333340
rect 82292 373072 82348 373184
rect 80836 255008 80892 333284
rect 82292 333228 82348 372624
rect 80948 333172 82348 333228
rect 82404 373072 82460 373184
rect 80948 255252 81004 333172
rect 82404 333116 82460 372624
rect 81060 333060 82460 333116
rect 82516 373072 82572 373184
rect 81060 255496 81116 333060
rect 82516 333004 82572 372624
rect 81172 332948 82572 333004
rect 82628 373072 82684 373184
rect 81172 255740 81228 332948
rect 82628 332892 82684 372624
rect 81284 332836 82684 332892
rect 82740 373072 82796 373184
rect 81284 255984 81340 332836
rect 82740 332780 82796 372624
rect 81396 332724 82796 332780
rect 82852 373072 82908 373184
rect 81396 258180 81452 332724
rect 82852 332668 82908 372624
rect 81508 332612 82908 332668
rect 82964 373072 83020 373184
rect 81508 258424 81564 332612
rect 82964 332556 83020 372624
rect 81620 332500 83020 332556
rect 83076 373072 83132 373184
rect 81620 258668 81676 332500
rect 83076 332444 83132 372624
rect 81732 332388 83132 332444
rect 83188 373072 83244 373184
rect 81732 258912 81788 332388
rect 83188 332332 83244 372624
rect 81844 332276 83244 332332
rect 83300 373072 83356 373184
rect 81844 259156 81900 332276
rect 83300 332220 83356 372624
rect 81956 332164 83356 332220
rect 83412 373072 83468 373184
rect 81956 259400 82012 332164
rect 83412 332108 83468 372624
rect 82068 332052 83468 332108
rect 83524 373072 83580 373184
rect 82068 259644 82124 332052
rect 83524 331996 83580 372624
rect 82180 331940 83580 331996
rect 83636 373072 83692 373184
rect 82180 259888 82236 331940
rect 83636 331884 83692 372624
rect 82292 331828 83692 331884
rect 83748 373072 83804 373184
rect 82292 260132 82348 331828
rect 83748 331772 83804 372624
rect 82404 331716 83804 331772
rect 83860 373072 83916 373184
rect 82404 260376 82460 331716
rect 83860 331660 83916 372624
rect 82516 331604 83916 331660
rect 83972 373072 84028 373184
rect 82516 260620 82572 331604
rect 83972 331548 84028 372624
rect 85428 373072 85484 373184
rect 84980 366150 85036 366240
rect 82628 331492 84028 331548
rect 84084 361270 84140 361310
rect 82628 266638 82684 331492
rect 84084 331212 84140 361214
rect 82740 331156 84140 331212
rect 84308 361026 84364 361066
rect 82740 286412 82796 331156
rect 84308 330988 84364 360970
rect 82740 286316 82796 286356
rect 82964 330932 84364 330988
rect 84532 360782 84588 360822
rect 82964 286300 83020 330932
rect 84532 330764 84588 360726
rect 82964 286204 83020 286244
rect 83188 330708 84588 330764
rect 84756 360538 84812 360578
rect 83188 286188 83244 330708
rect 84756 330540 84812 360482
rect 83188 286092 83244 286132
rect 83412 330484 84812 330540
rect 84980 348582 85036 366094
rect 85428 360294 85484 372624
rect 85428 360198 85484 360238
rect 85652 373072 85708 373184
rect 85652 360050 85708 372624
rect 85652 359940 85708 359994
rect 85876 373072 85932 373184
rect 85876 359806 85932 372624
rect 88424 371290 88480 371320
rect 87164 371038 87220 371098
rect 85876 359716 85932 359750
rect 86156 368834 86212 368874
rect 83412 286076 83468 330484
rect 84980 330316 85036 348526
rect 85358 348094 85414 348134
rect 83412 285964 83468 286020
rect 83636 330260 85036 330316
rect 85092 346630 85148 346668
rect 82628 266542 82684 266582
rect 82516 260524 82572 260564
rect 82404 260280 82460 260320
rect 82292 260036 82348 260076
rect 82180 259792 82236 259832
rect 82068 259548 82124 259588
rect 81956 259304 82012 259344
rect 81844 259060 81900 259100
rect 81732 258816 81788 258856
rect 81620 258572 81676 258612
rect 81508 258328 81564 258368
rect 81396 258084 81452 258124
rect 81284 255888 81340 255928
rect 81172 255644 81228 255684
rect 81060 255400 81116 255440
rect 80948 255156 81004 255196
rect 80836 254912 80892 254952
rect 80724 254668 80780 254708
rect 80612 254424 80668 254464
rect 80500 254180 80556 254220
rect 80388 253936 80444 253976
rect 80276 253692 80332 253732
rect 80164 253448 80220 253488
rect 80052 253204 80108 253244
rect 79940 252960 79996 253000
rect 79828 252716 79884 252756
rect 79716 252472 79772 252512
rect 79604 252228 79660 252268
rect 79492 251984 79548 252024
rect 79380 251740 79436 251780
rect 79268 251496 79324 251536
rect 79156 251252 79212 251292
rect 79044 251008 79100 251048
rect 78932 250764 78988 250804
rect 78820 250520 78876 250560
rect 78708 250276 78764 250316
rect 78596 249056 78652 249096
rect 78484 248812 78540 248852
rect 78372 248568 78428 248608
rect 78260 248324 78316 248364
rect 78148 248080 78204 248120
rect 78036 247836 78092 247876
rect 77924 247592 77980 247632
rect 77812 247348 77868 247388
rect 77700 247104 77756 247144
rect 77588 246860 77644 246900
rect 77476 246616 77532 246656
rect 77364 246372 77420 246412
rect 75012 246128 75068 246168
rect 74900 245884 74956 245924
rect 74788 245640 74844 245680
rect 74676 245396 74732 245436
rect 74452 239556 74508 239596
rect 73220 238868 83468 238924
rect 73108 238756 83356 238812
rect 72996 238644 83244 238700
rect 72884 238532 83132 238588
rect 72772 238420 83020 238476
rect 72660 238308 82908 238364
rect 72548 238196 82796 238252
rect 72436 238084 82684 238140
rect 72324 237972 82572 238028
rect 72212 237860 82460 237916
rect 72100 237748 82348 237804
rect 71988 237636 82236 237692
rect 71876 237524 82124 237580
rect 71764 237412 82012 237468
rect 71652 237300 81900 237356
rect 71540 237188 81788 237244
rect 71428 237076 81676 237132
rect 71316 236964 81564 237020
rect 71204 236852 81452 236908
rect 71092 236740 81340 236796
rect 70980 236628 81228 236684
rect 70868 236516 81116 236572
rect 70756 236404 81004 236460
rect 70644 236292 80892 236348
rect 70532 236180 80780 236236
rect 70420 236068 80668 236124
rect 70308 235956 80556 236012
rect 70196 235844 80444 235900
rect 70084 235732 80108 235788
rect 69972 235620 79996 235676
rect 69860 233940 70672 233996
rect 66276 233604 66780 233730
rect 66276 232596 66402 233604
rect 66654 232596 66780 233604
rect 66276 232470 66780 232596
rect 65306 232092 65347 232265
rect 65547 232092 66978 232265
rect 64917 231343 66977 231510
rect 64209 226767 64779 226800
rect 64209 225689 64234 226767
rect 64745 225689 64779 226767
rect 64209 225414 64779 225689
rect 64917 225382 65084 231343
rect 72324 229320 73710 229446
rect 72324 228690 72450 229320
rect 73584 228690 73710 229320
rect 72324 228564 73710 228690
rect 72828 209538 73710 209664
rect 72828 208656 72954 209538
rect 73584 208656 73710 209538
rect 72828 208530 73710 208656
rect 79254 207942 79758 208026
rect 35028 207508 36092 207564
rect 34895 206806 35247 206876
rect 34895 203662 34939 206806
rect 35194 203662 35247 206806
rect 34895 203610 35247 203662
rect 35495 190006 35847 190076
rect 35495 186862 35539 190006
rect 35794 186862 35847 190006
rect 35495 186810 35847 186862
rect 36036 174636 36092 207508
rect 79254 206980 79331 207942
rect 79685 206980 79758 207942
rect 79254 206892 79758 206980
rect 73444 206714 73500 206754
rect 37535 205873 39918 205885
rect 37535 205293 37590 205873
rect 38138 205293 39918 205873
rect 37535 205288 39918 205293
rect 73444 202104 73500 206658
rect 74116 206602 74172 206642
rect 73780 206000 73836 206046
rect 73780 203324 73836 205944
rect 73780 203240 73836 203268
rect 74116 202226 74172 206546
rect 74788 206490 74844 206530
rect 74306 205722 74654 205762
rect 74306 205038 74345 205722
rect 74614 205038 74654 205722
rect 74306 204996 74654 205038
rect 74788 202348 74844 206434
rect 75460 206378 75516 206418
rect 75124 206000 75180 206040
rect 75124 205258 75180 205944
rect 75124 205167 75180 205202
rect 75460 202470 75516 206322
rect 76132 206266 76188 206306
rect 75572 205370 75628 205412
rect 75572 203446 75628 205314
rect 75572 203347 75628 203390
rect 76132 202592 76188 206210
rect 76804 206154 76860 206194
rect 76804 202714 76860 206098
rect 77476 206042 77532 206082
rect 77364 205482 77420 205520
rect 77364 203568 77420 205426
rect 77364 203472 77420 203512
rect 77476 202836 77532 205986
rect 78148 205930 78204 205970
rect 78148 202958 78204 205874
rect 78820 205818 78876 205858
rect 78820 203080 78876 205762
rect 79492 205706 79548 205746
rect 79492 203202 79548 205650
rect 79492 203106 79548 203146
rect 78820 202984 78876 203024
rect 78148 202862 78204 202902
rect 77476 202756 77532 202780
rect 76804 202618 76860 202658
rect 76132 202496 76188 202536
rect 75460 202374 75516 202414
rect 74788 202252 74844 202292
rect 74116 202138 74172 202170
rect 73444 202008 73500 202048
rect 73080 200970 73836 201096
rect 70686 198940 71442 198976
rect 71587 198940 71903 200274
rect 71987 199900 72303 200274
rect 73080 199900 73206 200970
rect 71987 199710 73206 199900
rect 73710 199710 73836 200970
rect 71987 199584 73836 199710
rect 70686 198850 71903 198940
rect 64545 198350 64831 198372
rect 49770 197117 51912 197190
rect 49770 196869 49829 197117
rect 51830 196869 51912 197117
rect 49770 196812 51912 196869
rect 49840 196492 50440 196812
rect 37707 195078 39954 195086
rect 37707 194653 37740 195078
rect 38303 194653 39954 195078
rect 37707 194651 39954 194653
rect 64545 187864 64831 198151
rect 70686 198094 70812 198850
rect 71316 198624 71903 198850
rect 71316 198094 71442 198624
rect 70686 197968 71442 198094
rect 65443 197670 65722 197766
rect 65443 191212 65722 197377
rect 68922 193032 69678 193158
rect 68922 192402 69048 193032
rect 69552 192402 69678 193032
rect 68922 192276 69678 192402
rect 79940 191772 79996 235620
rect 69748 191716 79996 191772
rect 65443 191018 67079 191212
rect 69748 190932 69804 191716
rect 80052 191660 80108 235732
rect 80164 205594 80220 205634
rect 80164 203690 80220 205538
rect 80164 203604 80220 203634
rect 70756 191604 80108 191660
rect 70756 190932 70812 191604
rect 66024 190008 66906 190134
rect 66024 189252 66150 190008
rect 66780 189252 66906 190008
rect 66024 189126 66906 189252
rect 64545 187617 64831 187664
rect 64921 188434 67095 188574
rect 64228 184338 64780 184386
rect 64228 182952 64260 184338
rect 64764 182952 64780 184338
rect 64228 182619 64780 182952
rect 64180 182574 64780 182619
rect 64921 182595 65061 188434
rect 66770 185968 67122 185991
rect 66770 185801 66801 185968
rect 67096 185801 67122 185968
rect 66770 185782 67122 185801
rect 36036 174580 37212 174636
rect 36095 173206 36447 173276
rect 36095 170062 36139 173206
rect 36394 170062 36447 173206
rect 36095 170010 36447 170062
rect 36695 156406 37047 156476
rect 36695 153262 36739 156406
rect 36994 153262 37047 156406
rect 36695 153210 37047 153262
rect 32998 146076 33054 146116
rect 32550 119202 32606 122368
rect 32550 118836 32606 118958
rect 32802 145816 32858 145856
rect 32802 143388 32858 145760
rect 32998 143612 33054 146020
rect 37156 146076 37212 174580
rect 73206 167202 74214 167328
rect 73206 166446 73332 167202
rect 74088 166446 74214 167202
rect 73206 166320 74214 166446
rect 79380 165312 80010 165438
rect 79380 164178 79506 165312
rect 79884 164178 80010 165312
rect 79380 164052 80010 164178
rect 73444 163892 73500 163932
rect 37535 163073 39920 163085
rect 37535 162493 37590 163073
rect 38138 162493 39920 163073
rect 37535 162488 39920 162493
rect 73444 159282 73500 163836
rect 80388 163892 80444 235844
rect 74116 163780 74172 163820
rect 80388 163796 80444 163836
rect 73780 162436 73836 162474
rect 73780 160502 73836 162380
rect 73780 160418 73836 160446
rect 74116 159404 74172 163724
rect 80500 163780 80556 235956
rect 74788 163668 74844 163708
rect 80500 163684 80556 163724
rect 74788 159526 74844 163612
rect 80612 163668 80668 236068
rect 75460 163556 75516 163596
rect 80612 163572 80668 163612
rect 75460 159648 75516 163500
rect 80724 163556 80780 236180
rect 76132 163444 76188 163484
rect 80724 163460 80780 163500
rect 75572 162548 75628 162586
rect 75572 160624 75628 162492
rect 75572 160525 75628 160568
rect 76132 159770 76188 163388
rect 80836 163444 80892 236292
rect 76804 163332 76860 163372
rect 80836 163348 80892 163388
rect 76804 159892 76860 163276
rect 80948 163332 81004 236404
rect 77476 163220 77532 163260
rect 80948 163236 81004 163276
rect 77364 162660 77420 162692
rect 77364 160746 77420 162604
rect 77364 160650 77420 160690
rect 77476 160014 77532 163164
rect 81060 163220 81116 236516
rect 78148 163108 78204 163148
rect 81060 163124 81116 163164
rect 78148 160136 78204 163052
rect 81172 163108 81228 236628
rect 78820 162996 78876 163036
rect 81172 163012 81228 163052
rect 78820 160258 78876 162940
rect 81284 162996 81340 236740
rect 79492 162884 79548 162924
rect 81284 162900 81340 162940
rect 79492 160380 79548 162828
rect 81396 162884 81452 236852
rect 80164 162772 80220 162812
rect 81396 162788 81452 162828
rect 80164 160868 80220 162716
rect 81508 162772 81564 236964
rect 81508 162676 81564 162716
rect 81620 162660 81676 237076
rect 81620 162564 81676 162604
rect 81732 162548 81788 237188
rect 81732 162452 81788 162492
rect 81844 162436 81900 237300
rect 81956 206714 82012 237412
rect 81956 206618 82012 206658
rect 82068 206602 82124 237524
rect 82068 206506 82124 206546
rect 82180 206490 82236 237636
rect 82180 206394 82236 206434
rect 82292 206378 82348 237748
rect 82292 206282 82348 206322
rect 82404 206266 82460 237860
rect 82404 206170 82460 206210
rect 82516 206154 82572 237972
rect 82516 206058 82572 206098
rect 82628 206042 82684 238084
rect 82628 205946 82684 205986
rect 82740 205930 82796 238196
rect 82740 205834 82796 205874
rect 82852 205818 82908 238308
rect 82852 205722 82908 205762
rect 82964 205706 83020 238420
rect 82964 205610 83020 205650
rect 83076 205594 83132 238532
rect 83076 205498 83132 205538
rect 83188 205482 83244 238644
rect 83188 205386 83244 205426
rect 83300 205370 83356 238756
rect 83300 205274 83356 205314
rect 83412 205258 83468 238868
rect 83412 205162 83468 205202
rect 81844 162340 81900 162380
rect 80766 162036 81648 162162
rect 80766 161532 80892 162036
rect 81522 161532 81648 162036
rect 80766 161406 81648 161532
rect 80164 160772 80220 160812
rect 79492 160284 79548 160324
rect 78820 160162 78876 160202
rect 78148 160040 78204 160080
rect 77476 159920 77532 159958
rect 76804 159796 76860 159836
rect 76132 159674 76188 159714
rect 75460 159552 75516 159592
rect 74788 159430 74844 159470
rect 74116 159296 74172 159348
rect 73444 159186 73500 159226
rect 70880 156878 71196 156880
rect 71588 156878 71904 157448
rect 70878 156752 71904 156878
rect 71988 156870 72304 157448
rect 70878 156500 70964 156752
rect 71720 156500 71904 156752
rect 70878 156376 71904 156500
rect 71986 156744 72954 156870
rect 71986 156492 72072 156744
rect 72828 156492 72954 156744
rect 70878 156374 71108 156376
rect 70880 156373 71108 156374
rect 71986 156366 72954 156492
rect 71988 156365 72304 156366
rect 61684 155596 61740 155606
rect 60004 155456 60060 155496
rect 51282 153468 52920 153594
rect 51282 152838 51408 153468
rect 52794 152838 52920 153468
rect 51282 152712 52920 152838
rect 52164 148371 52220 148405
rect 37156 146010 37212 146020
rect 47236 145964 47292 146188
rect 47236 145796 47292 145908
rect 52164 145824 52220 148226
rect 52724 148370 52780 148405
rect 52500 146848 52556 146890
rect 52500 146636 52556 146702
rect 52500 145824 52556 146580
rect 52724 145824 52780 148226
rect 53284 148370 53340 148405
rect 53060 146848 53116 146890
rect 53060 146412 53116 146702
rect 53060 145824 53116 146356
rect 53284 145824 53340 148226
rect 53844 148370 53900 148405
rect 53620 146848 53676 146880
rect 53620 146188 53676 146702
rect 53620 145824 53676 146132
rect 53844 145824 53900 148217
rect 54180 146848 54236 146888
rect 54180 145964 54236 146702
rect 54180 145824 54236 145908
rect 55524 146188 55580 146832
rect 55524 145796 55580 146132
rect 56644 146412 56700 146832
rect 56644 145796 56700 146356
rect 56868 146636 56924 146832
rect 56868 145796 56924 146580
rect 32998 143492 33054 143556
rect 32802 119202 32858 143332
rect 32802 118836 32858 118958
rect 33054 143164 33110 143204
rect 33054 119202 33110 143108
rect 33054 118836 33110 118958
rect 33306 142940 33362 142980
rect 33306 119202 33362 142884
rect 33306 118836 33362 118958
rect 33558 142716 33614 142756
rect 33558 119202 33614 142660
rect 33558 118836 33614 118958
rect 33810 142492 33866 142532
rect 33810 119202 33866 142436
rect 58548 140028 58604 140068
rect 58324 137340 58380 137380
rect 44324 122668 44380 124792
rect 48916 122892 48972 124792
rect 51828 123116 51884 124792
rect 52052 123340 52108 124792
rect 52276 123564 52332 124792
rect 52500 123788 52556 124792
rect 52500 123536 52556 123732
rect 52724 124012 52780 124792
rect 52724 123536 52780 123956
rect 53284 124236 53340 124792
rect 53284 123536 53340 124180
rect 56308 124460 56364 124792
rect 56308 123536 56364 124404
rect 52276 123468 52332 123508
rect 52052 123244 52108 123284
rect 51828 123020 51884 123060
rect 48916 122796 48972 122836
rect 44324 122572 44380 122612
rect 39360 121548 39428 121588
rect 39232 121324 39300 121364
rect 39104 121100 39172 121140
rect 33810 118836 33866 118958
rect 38976 120876 39044 120916
rect 32200 116175 34542 117908
rect 32200 116046 37855 116175
rect 32200 114912 34650 116046
rect 35406 114912 37855 116046
rect 32200 114788 37855 114912
rect 32200 109085 34542 114788
rect 32200 101246 34333 109085
rect 34506 101246 34542 109085
rect 37548 109620 38682 109746
rect 37548 108612 37674 109620
rect 38556 108612 38682 109620
rect 37548 108486 38682 108612
rect 32200 76798 34542 101246
rect 35188 107984 37870 108040
rect 38167 107984 38192 108040
rect 35188 95584 35244 107984
rect 35188 95468 35244 95508
rect 35524 107648 37870 107704
rect 38167 107648 38192 107704
rect 35524 78178 35580 107648
rect 38976 105964 39044 120820
rect 39104 105964 39172 121044
rect 39232 105964 39300 121268
rect 39360 105964 39428 121492
rect 58324 108040 58380 137284
rect 58548 130995 58604 139972
rect 58548 130947 58621 130995
rect 58548 130697 58556 130947
rect 58620 130697 58621 130947
rect 60004 130878 60060 155400
rect 61334 144966 61390 145086
rect 61334 143866 61390 144890
rect 61684 145040 61740 155540
rect 61684 144676 61740 144816
rect 61796 155334 61852 155374
rect 61334 143800 61390 143810
rect 61796 136556 61852 155278
rect 62356 155212 62412 155252
rect 62356 145040 62412 155156
rect 61908 144956 61964 145040
rect 61908 139132 61964 144900
rect 62356 144676 62412 144816
rect 62468 155090 62524 155130
rect 61908 139036 61964 139076
rect 62468 136556 62524 155034
rect 63028 154968 63084 155008
rect 63028 145040 63084 154912
rect 62580 144956 62636 145040
rect 62580 138908 62636 144900
rect 63028 144676 63084 144816
rect 63140 154846 63196 154886
rect 62580 138812 62636 138852
rect 61684 136500 61852 136556
rect 62244 136500 62524 136556
rect 63140 136546 63196 154790
rect 63700 154724 63756 154764
rect 63700 145040 63756 154668
rect 63252 144956 63308 145040
rect 63252 138684 63308 144900
rect 63700 144676 63756 144816
rect 63812 154602 63868 154642
rect 63252 138588 63308 138628
rect 63812 136668 63868 154546
rect 64372 154480 64428 154520
rect 64372 145040 64428 154424
rect 63924 144956 63980 145040
rect 63924 138460 63980 144900
rect 64372 144676 64428 144816
rect 64484 154358 64540 154398
rect 63924 138364 63980 138404
rect 60858 135828 61488 135954
rect 60858 133560 60984 135828
rect 61362 133560 61488 135828
rect 61684 134428 61740 136500
rect 62244 135546 62300 136500
rect 61908 135436 61964 135476
rect 61908 134652 61964 135380
rect 62916 136490 63196 136546
rect 63588 136612 63868 136668
rect 62916 135546 62972 136490
rect 62244 135156 62300 135268
rect 62580 135436 62636 135476
rect 62580 134988 62636 135380
rect 63588 135546 63644 136612
rect 64484 136556 64540 154302
rect 65044 154236 65100 154276
rect 65044 145040 65100 154180
rect 64596 144956 64652 145040
rect 64596 138236 64652 144900
rect 65044 144676 65100 144816
rect 65156 154114 65212 154154
rect 64596 138140 64652 138180
rect 65156 136556 65212 154058
rect 65716 153992 65772 154032
rect 65716 145040 65772 153936
rect 65268 144956 65324 145040
rect 65268 138012 65324 144900
rect 65716 144676 65772 144816
rect 65828 153870 65884 153910
rect 65268 137916 65324 137956
rect 65828 136556 65884 153814
rect 66388 153748 66444 153788
rect 66388 145040 66444 153692
rect 65940 144956 65996 145040
rect 65940 137788 65996 144900
rect 66388 144676 66444 144816
rect 66500 153626 66556 153666
rect 65940 137692 65996 137732
rect 66500 136556 66556 153570
rect 67060 153504 67116 153544
rect 67060 145040 67116 153448
rect 66612 144956 66668 145040
rect 66612 137564 66668 144900
rect 67060 144676 67116 144816
rect 67172 153382 67228 153422
rect 66612 137468 66668 137508
rect 67172 136556 67228 153326
rect 67732 153260 67788 153300
rect 67732 145040 67788 153204
rect 67284 144956 67340 145040
rect 67284 142716 67340 144900
rect 67732 144676 67788 144816
rect 67844 153138 67900 153178
rect 67284 142620 67340 142660
rect 67844 136892 67900 153082
rect 68404 152894 68460 152934
rect 68404 145040 68460 152838
rect 68850 152772 68910 152812
rect 67956 144956 68012 145040
rect 67956 142492 68012 144900
rect 68404 144676 68460 144816
rect 68628 144956 68684 145040
rect 67956 142396 68012 142436
rect 68628 142268 68684 144900
rect 68628 142172 68684 142212
rect 68850 139134 68910 152716
rect 69076 152650 69132 152690
rect 69076 145040 69132 152594
rect 69636 152528 69692 152568
rect 69076 144676 69132 144816
rect 69300 144956 69356 145040
rect 69300 142044 69356 144900
rect 69300 141948 69356 141988
rect 62916 135156 62972 135268
rect 63252 135436 63308 135476
rect 62580 134932 62748 134988
rect 61908 134596 62188 134652
rect 61684 134372 61852 134428
rect 60858 133434 61488 133560
rect 58548 130650 58621 130697
rect 59960 130853 60060 130878
rect 60016 130683 60060 130853
rect 59960 130656 60060 130683
rect 58548 130564 58604 130650
rect 60004 130637 60060 130656
rect 60340 130930 60396 131040
rect 60340 130906 60409 130930
rect 60340 130736 60353 130906
rect 61796 130875 61852 134372
rect 62132 133411 62188 134596
rect 62132 133229 62188 133262
rect 62692 133411 62748 134932
rect 62692 133229 62748 133262
rect 63252 133411 63308 135380
rect 64260 136500 64540 136556
rect 64932 136500 65212 136556
rect 65604 136500 65884 136556
rect 66276 136500 66556 136556
rect 66948 136500 67228 136556
rect 67620 136836 67900 136892
rect 68628 139074 68910 139134
rect 64260 135546 64316 136500
rect 63588 135156 63644 135268
rect 63924 135436 63980 135476
rect 63924 134988 63980 135380
rect 64932 135546 64988 136500
rect 64260 135156 64316 135268
rect 64596 135436 64652 135476
rect 64596 134988 64652 135380
rect 65604 135546 65660 136500
rect 64932 135156 64988 135268
rect 65268 135436 65324 135476
rect 63252 133229 63308 133262
rect 63812 134932 63980 134988
rect 64372 134932 64652 134988
rect 63812 133411 63868 134932
rect 63812 133229 63868 133262
rect 64372 133416 64428 134932
rect 65268 134764 65324 135380
rect 66276 135546 66332 136500
rect 65604 135156 65660 135268
rect 65940 135436 65996 135476
rect 64372 133229 64428 133257
rect 64932 134708 65324 134764
rect 64932 133416 64988 134708
rect 65940 134540 65996 135380
rect 66948 135546 67004 136500
rect 66276 135156 66332 135268
rect 66612 135436 66668 135476
rect 64932 133229 64988 133257
rect 65492 134484 65996 134540
rect 65492 133416 65548 134484
rect 66612 134316 66668 135380
rect 67620 135546 67676 136836
rect 66948 135156 67004 135268
rect 67284 135436 67340 135520
rect 67284 134540 67340 135380
rect 68292 135546 68348 136668
rect 67620 135156 67676 135268
rect 67956 135436 68012 135520
rect 67284 134484 67452 134540
rect 65492 133229 65548 133257
rect 66052 134260 66668 134316
rect 66052 133416 66108 134260
rect 66052 133229 66108 133257
rect 66612 133416 66668 133504
rect 66612 131964 66668 133257
rect 62622 131292 65772 131418
rect 62622 131040 62748 131292
rect 65646 131040 65772 131292
rect 62622 130914 65772 131040
rect 60340 130708 60409 130736
rect 61755 130853 61852 130875
rect 59850 130511 60099 130525
rect 59850 130503 59875 130511
rect 60078 130503 60099 130511
rect 59760 130447 59780 130503
rect 60083 130447 60099 130503
rect 59850 130057 59875 130447
rect 60078 130057 60099 130447
rect 59850 130032 60099 130057
rect 60340 128044 60396 130708
rect 61811 130683 61852 130853
rect 61755 130658 61852 130683
rect 61796 130630 61852 130658
rect 61562 130445 61577 130502
rect 61880 130445 61902 130502
rect 61611 130051 61634 130445
rect 61874 130051 61902 130445
rect 61611 130030 61902 130051
rect 62622 130410 65772 130536
rect 62622 130158 62748 130410
rect 65646 130158 65772 130410
rect 62622 130032 65772 130158
rect 60340 127904 60396 127988
rect 59724 127638 60228 127764
rect 59724 127386 59850 127638
rect 60102 127386 60228 127638
rect 59114 127246 59194 127279
rect 59724 127260 60228 127386
rect 59114 127082 59115 127246
rect 59193 127082 59194 127246
rect 59114 124684 59194 127082
rect 60984 127008 61992 127134
rect 60984 126630 61110 127008
rect 61866 126630 61992 127008
rect 60984 126504 61992 126630
rect 59114 124616 59194 124628
rect 66612 124908 66668 131908
rect 67172 133416 67228 133504
rect 67172 131964 67228 133257
rect 67172 131898 67228 131908
rect 67396 126252 67452 134484
rect 67956 134316 68012 135380
rect 68292 135156 68348 135268
rect 68628 135546 68684 139074
rect 69636 135546 69692 152472
rect 69748 152406 69804 152446
rect 69748 145040 69804 152350
rect 70308 152284 70364 152324
rect 69748 144676 69804 144816
rect 69972 144956 70028 145040
rect 69972 141820 70028 144900
rect 69972 141724 70028 141764
rect 68628 135156 68684 135268
rect 68964 135436 69020 135520
rect 67732 134260 68012 134316
rect 67732 133416 67788 134260
rect 67732 133084 67788 133257
rect 68292 133416 68348 133504
rect 68292 133084 68348 133257
rect 67732 133028 68348 133084
rect 68852 133416 68908 133504
rect 67732 131964 67788 133028
rect 67732 131898 67788 131908
rect 68852 131964 68908 133257
rect 68852 131898 68908 131908
rect 68964 130633 69020 135380
rect 68964 128940 69020 130577
rect 68964 128844 69020 128884
rect 69188 135436 69244 135520
rect 69188 128268 69244 135380
rect 70308 135546 70364 152228
rect 70420 152162 70476 152202
rect 70420 145040 70476 152106
rect 70980 152040 71036 152080
rect 70420 144676 70476 144816
rect 70644 144956 70700 145040
rect 70644 141596 70700 144900
rect 70644 141500 70700 141540
rect 69636 135156 69692 135268
rect 69860 135436 69916 135520
rect 69412 133416 69468 133504
rect 69412 131964 69468 133257
rect 69412 131898 69468 131908
rect 69860 129836 69916 135380
rect 70532 136332 70588 136416
rect 70532 135436 70588 136276
rect 70532 135296 70588 135380
rect 70980 135546 71036 151984
rect 71092 151918 71148 151958
rect 71092 145040 71148 151862
rect 71652 151796 71708 151836
rect 71092 144676 71148 144816
rect 71316 144956 71372 145040
rect 71316 141372 71372 144900
rect 71316 141276 71372 141316
rect 70308 135156 70364 135268
rect 71204 136108 71260 136192
rect 71204 135436 71260 136052
rect 71204 135296 71260 135380
rect 71652 135546 71708 151740
rect 71764 151674 71820 151714
rect 71764 145040 71820 151618
rect 72324 151552 72380 151592
rect 71764 144676 71820 144816
rect 71988 144956 72044 145040
rect 71988 141148 72044 144900
rect 71988 141052 72044 141092
rect 69972 133416 70028 133504
rect 69972 131964 70028 133257
rect 69972 131898 70028 131908
rect 70532 133416 70588 133504
rect 70532 131964 70588 133257
rect 70532 131898 70588 131908
rect 69860 129740 69916 129780
rect 69188 128172 69244 128212
rect 67396 126156 67452 126196
rect 66612 122424 66668 124852
rect 66612 122328 66668 122368
rect 70550 121772 70606 121782
rect 63513 111591 65199 111650
rect 63513 111371 63569 111591
rect 65143 111556 65199 111591
rect 63513 111250 63569 111275
rect 63875 111474 63931 111488
rect 58324 107940 58380 107984
rect 59000 110110 59056 110158
rect 39560 106605 39628 106627
rect 39560 105964 39628 106453
rect 41220 106310 41288 106336
rect 41220 105970 41288 106254
rect 59000 106310 59056 110054
rect 61455 108515 61468 108571
rect 61636 108515 61653 108571
rect 63875 108559 63931 111368
rect 64889 111352 64945 111369
rect 65143 111256 65199 111308
rect 66033 111591 67719 111650
rect 66033 111371 66089 111591
rect 67663 111556 67719 111591
rect 66033 111250 66089 111275
rect 66395 111474 66451 111497
rect 64889 111131 64945 111196
rect 66395 111131 66451 111368
rect 64889 111075 66451 111131
rect 67409 111352 67465 111369
rect 67663 111256 67719 111308
rect 68553 111591 70239 111650
rect 68553 111371 68609 111591
rect 70183 111556 70239 111591
rect 68553 111250 68609 111275
rect 68915 111474 68971 111497
rect 67409 111131 67465 111196
rect 68915 111131 68971 111368
rect 67409 111075 68971 111131
rect 69929 111352 69985 111369
rect 70183 111256 70239 111308
rect 69929 111131 69985 111196
rect 70550 111131 70606 121716
rect 69929 111075 70606 111131
rect 70980 110110 71036 135268
rect 70980 110004 71036 110054
rect 72324 135546 72380 151496
rect 72436 151430 72492 151470
rect 72436 145040 72492 151374
rect 72996 151308 73052 151348
rect 72436 144676 72492 144816
rect 72660 144956 72716 145040
rect 72660 140924 72716 144900
rect 72660 140828 72716 140868
rect 66780 109116 67662 109242
rect 66780 108738 66906 109116
rect 67536 108738 67662 109116
rect 66780 108612 67662 108738
rect 68152 108581 68212 108609
rect 61486 107704 61546 108515
rect 63827 108503 63850 108559
rect 64165 108503 64190 108559
rect 61486 107628 61546 107648
rect 59472 107352 60732 107478
rect 59472 106974 59598 107352
rect 60606 106974 60732 107352
rect 59472 106848 60732 106974
rect 63875 106886 63931 108503
rect 70980 108500 71008 108556
rect 71450 108500 71478 108556
rect 65772 107604 66654 107730
rect 65772 107226 65898 107604
rect 66528 107226 66654 107604
rect 68152 107646 68212 108469
rect 68152 107590 68592 107646
rect 65772 107100 66654 107226
rect 63875 106830 68212 106886
rect 59000 106200 59056 106254
rect 62364 106198 62384 106254
rect 62658 106198 62674 106254
rect 62486 105963 62546 106198
rect 68152 105957 68212 106830
rect 68536 106254 68592 107590
rect 71652 106304 71708 135268
rect 71876 135436 71932 135520
rect 71876 131628 71932 135380
rect 72548 137340 72604 137424
rect 72548 135436 72604 137284
rect 72548 135296 72604 135380
rect 72996 135546 73052 151252
rect 73108 151186 73164 151226
rect 73108 145040 73164 151130
rect 73668 151064 73724 151104
rect 73108 144676 73164 144816
rect 73332 144956 73388 145040
rect 73332 140700 73388 144900
rect 73332 140604 73388 140644
rect 72324 133284 72380 135268
rect 73220 137116 73276 137200
rect 73220 135436 73276 137060
rect 73220 135296 73276 135380
rect 73668 135546 73724 151008
rect 73780 150942 73836 150982
rect 73780 145040 73836 150886
rect 74340 150820 74396 150860
rect 73780 144676 73836 144816
rect 74004 144956 74060 145040
rect 74004 140476 74060 144900
rect 74004 140380 74060 140420
rect 72996 135156 73052 135268
rect 74340 135546 74396 150764
rect 74452 150698 74508 150738
rect 74452 145040 74508 150642
rect 75012 150576 75068 150616
rect 74452 144676 74508 144816
rect 74676 144956 74732 145040
rect 74676 140252 74732 144900
rect 74676 140156 74732 140196
rect 73668 135156 73724 135268
rect 73892 135436 73948 135520
rect 72324 133228 73528 133284
rect 72188 132804 73196 132930
rect 72188 132174 72314 132804
rect 73070 132174 73196 132804
rect 72188 132048 73196 132174
rect 71876 131532 71932 131572
rect 73472 106746 73528 133228
rect 73892 124460 73948 135380
rect 73892 124364 73948 124404
rect 75012 135546 75068 150520
rect 75124 150454 75180 150494
rect 75124 145040 75180 150398
rect 75684 150332 75740 150372
rect 75124 144676 75180 144816
rect 75348 144956 75404 145040
rect 75348 143612 75404 144900
rect 75348 143516 75404 143556
rect 74340 121548 74396 135268
rect 74564 135436 74620 135520
rect 74564 124236 74620 135380
rect 74564 124140 74620 124180
rect 75684 135546 75740 150276
rect 75796 150210 75852 150250
rect 75796 145040 75852 150154
rect 76356 150088 76412 150128
rect 75796 144676 75852 144816
rect 76020 144956 76076 145040
rect 76020 143388 76076 144900
rect 76020 143292 76076 143332
rect 74340 121482 74396 121492
rect 75012 121324 75068 135268
rect 75236 135436 75292 135520
rect 75236 124012 75292 135380
rect 75236 123916 75292 123956
rect 76356 135546 76412 150032
rect 76468 149966 76524 150006
rect 76468 145040 76524 149910
rect 77028 149844 77084 149884
rect 76468 144676 76524 144816
rect 76692 144956 76748 145040
rect 76692 143164 76748 144900
rect 76692 143068 76748 143108
rect 75012 121258 75068 121268
rect 75684 121100 75740 135268
rect 75908 135436 75964 135520
rect 75908 123788 75964 135380
rect 75908 123692 75964 123732
rect 77028 135546 77084 149788
rect 77140 149722 77196 149762
rect 77140 145040 77196 149666
rect 77812 149600 77868 149640
rect 77812 145040 77868 149544
rect 78484 149478 78540 149518
rect 78484 145040 78540 149422
rect 79156 149356 79212 149396
rect 79156 145040 79212 149300
rect 79828 149234 79884 149274
rect 79828 145040 79884 149178
rect 77140 144676 77196 144816
rect 77364 144956 77420 145040
rect 77364 142940 77420 144900
rect 77812 144676 77868 144816
rect 78036 144956 78092 145040
rect 77364 142844 77420 142884
rect 78036 139804 78092 144900
rect 78484 144676 78540 144816
rect 78708 144956 78764 145040
rect 78036 139708 78092 139748
rect 78708 139580 78764 144900
rect 79156 144676 79212 144816
rect 79380 144956 79436 145040
rect 78708 139484 78764 139524
rect 79380 139356 79436 144900
rect 79828 144676 79884 144816
rect 80500 148136 80556 148176
rect 79380 139260 79436 139300
rect 75684 121034 75740 121044
rect 76356 120876 76412 135268
rect 76580 135436 76636 135520
rect 76580 122668 76636 135380
rect 77700 135546 77756 135632
rect 77028 135156 77084 135268
rect 77252 135436 77308 135520
rect 77252 123564 77308 135380
rect 77252 123468 77308 123508
rect 78372 135546 78428 135632
rect 76580 122572 76636 122612
rect 77700 121996 77756 135268
rect 77924 135436 77980 135520
rect 77924 123340 77980 135380
rect 77924 123244 77980 123284
rect 79044 135546 79100 135632
rect 78372 122220 78428 135268
rect 78596 135436 78652 135520
rect 78596 123116 78652 135380
rect 78596 123020 78652 123060
rect 79716 135546 79772 135632
rect 79044 122444 79100 135268
rect 79268 135436 79324 135520
rect 79268 122892 79324 135380
rect 79268 122796 79324 122836
rect 79716 122668 79772 135268
rect 79716 122572 79772 122612
rect 79044 122348 79100 122388
rect 78372 122124 78428 122164
rect 77700 121900 77756 121940
rect 80500 121772 80556 148080
rect 80500 121676 80556 121716
rect 80836 147892 80892 147932
rect 76356 120810 76412 120820
rect 80836 108556 80892 147836
rect 81144 146412 81774 146538
rect 81144 142380 81270 146412
rect 81648 142380 81774 146412
rect 82432 144978 83216 145040
rect 82432 144633 82494 144978
rect 83152 144633 83216 144978
rect 82432 144592 83216 144633
rect 81144 136458 81774 142380
rect 83636 137368 83692 330260
rect 85092 330204 85148 346574
rect 83748 330148 85148 330204
rect 83748 155596 83804 330148
rect 85358 329938 85414 348038
rect 84014 329882 85414 329938
rect 83748 155530 83804 155540
rect 83888 197342 83944 197361
rect 83888 155456 83944 197286
rect 83888 155334 83944 155400
rect 84014 155334 84070 329882
rect 86030 316618 86086 316658
rect 85778 316374 85834 316414
rect 85526 316130 85582 316170
rect 85274 315886 85330 315926
rect 85022 315642 85078 315682
rect 84770 315398 84826 315438
rect 84518 315154 84574 315194
rect 84266 314910 84322 314950
rect 84014 155238 84070 155278
rect 84140 305638 84196 305678
rect 84140 155212 84196 305582
rect 84140 155116 84196 155156
rect 84266 155090 84322 314854
rect 84266 154994 84322 155034
rect 84392 313202 84448 313242
rect 84392 154968 84448 313146
rect 84392 154872 84448 154912
rect 84518 154846 84574 315098
rect 84518 154750 84574 154790
rect 84644 313446 84700 313486
rect 84644 154724 84700 313390
rect 84644 154628 84700 154668
rect 84770 154602 84826 315342
rect 84770 154506 84826 154546
rect 84896 313690 84952 313730
rect 84896 154480 84952 313634
rect 84896 154384 84952 154424
rect 85022 154358 85078 315586
rect 85022 154262 85078 154302
rect 85148 313934 85204 313974
rect 85148 154236 85204 313878
rect 85148 154140 85204 154180
rect 85274 154114 85330 315830
rect 85274 154018 85330 154058
rect 85400 314178 85456 314218
rect 85400 153992 85456 314122
rect 85400 153896 85456 153936
rect 85526 153870 85582 316074
rect 85526 153774 85582 153814
rect 85652 314422 85708 314462
rect 85652 153748 85708 314366
rect 85652 153652 85708 153692
rect 85778 153626 85834 316318
rect 85778 153530 85834 153570
rect 85904 314666 85960 314706
rect 85904 153504 85960 314610
rect 85904 153408 85960 153448
rect 86030 153382 86086 316562
rect 86030 153286 86086 153326
rect 86156 153260 86212 368778
rect 86534 368590 86590 368630
rect 86408 348338 86464 348367
rect 86156 153164 86212 153204
rect 86282 317838 86338 317878
rect 86282 153138 86338 317782
rect 86282 153056 86338 153082
rect 86156 153016 86212 153056
rect 84870 147644 84926 147666
rect 84422 146972 84478 146995
rect 84422 145361 84478 146916
rect 84870 145361 84926 147588
rect 86156 147644 86212 152960
rect 86408 148639 86464 348282
rect 86534 152894 86590 368534
rect 86786 368346 86842 368386
rect 86534 152798 86590 152838
rect 86660 347606 86716 347630
rect 86660 152772 86716 347550
rect 86660 152678 86716 152716
rect 86786 152650 86842 368290
rect 87038 368102 87094 368142
rect 86786 152554 86842 152594
rect 86912 348826 86968 348866
rect 86912 152528 86968 348770
rect 86912 152432 86968 152472
rect 87038 152406 87094 368046
rect 87164 153016 87220 370982
rect 87164 152920 87220 152960
rect 87290 367858 87346 367898
rect 87038 152310 87094 152350
rect 87164 152284 87220 152324
rect 86408 148583 87024 148639
rect 86156 147578 86212 147588
rect 85990 147420 86046 147447
rect 84646 145226 84663 145302
rect 84797 145226 84814 145302
rect 84422 145152 84478 145174
rect 84706 145034 84762 145226
rect 85318 146972 85374 146992
rect 85318 145361 85374 146916
rect 85094 145226 85111 145302
rect 85245 145226 85262 145302
rect 84870 145152 84926 145174
rect 85154 145034 85210 145226
rect 85990 145353 86046 147364
rect 85542 145226 85559 145302
rect 85693 145226 85710 145302
rect 85318 145152 85374 145174
rect 85652 145034 85708 145226
rect 86662 147196 86718 147228
rect 86662 145353 86718 147140
rect 86214 145226 86231 145302
rect 86365 145226 86382 145302
rect 85990 145144 86046 145166
rect 86243 145034 86299 145226
rect 86662 145144 86718 145166
rect 84706 144978 86338 145034
rect 83636 137263 83692 137312
rect 81144 134946 81270 136458
rect 81648 134946 81774 136458
rect 81144 134820 81774 134946
rect 86282 130633 86338 144978
rect 86968 137766 87024 148583
rect 87164 147648 87220 152228
rect 87290 152162 87346 367802
rect 87542 367614 87598 367654
rect 87290 152066 87346 152106
rect 87416 347118 87472 347158
rect 87416 152040 87472 347062
rect 87416 151944 87472 151984
rect 87542 151918 87598 367558
rect 87794 367370 87850 367410
rect 87542 151822 87598 151862
rect 87668 347362 87724 347402
rect 87668 151796 87724 347306
rect 87668 151700 87724 151740
rect 87794 151674 87850 367314
rect 88046 367126 88102 367166
rect 87794 151578 87850 151618
rect 87920 346874 87976 346914
rect 87920 151552 87976 346818
rect 87920 151456 87976 151496
rect 88046 151430 88102 367070
rect 88298 366882 88354 366922
rect 88046 151334 88102 151374
rect 88172 347850 88228 347890
rect 88172 151308 88228 347794
rect 88172 151212 88228 151252
rect 88298 151186 88354 366826
rect 88298 151104 88354 151130
rect 88046 151064 88102 151104
rect 87154 147592 87164 147648
rect 87220 147592 87230 147648
rect 88046 146682 88102 151008
rect 88424 147420 88480 371234
rect 88676 370298 88732 370338
rect 88550 366638 88606 366678
rect 88550 150942 88606 366582
rect 88550 150846 88606 150886
rect 88676 150820 88732 370242
rect 88928 370054 88984 370094
rect 88676 150724 88732 150764
rect 88802 366394 88858 366434
rect 88802 150698 88858 366338
rect 88802 150602 88858 150642
rect 88928 150576 88984 369998
rect 89180 369810 89236 369850
rect 88928 150480 88984 150520
rect 89054 366150 89110 366190
rect 89054 150454 89110 366094
rect 89054 150358 89110 150398
rect 89180 150332 89236 369754
rect 89432 369566 89488 369606
rect 89180 150236 89236 150276
rect 89306 317594 89362 317634
rect 89306 150210 89362 317538
rect 89306 150114 89362 150154
rect 89432 150088 89488 369510
rect 90468 365174 90524 365214
rect 89798 356090 89824 356146
rect 90170 356090 90192 356146
rect 89798 355846 89824 355902
rect 90170 355846 90192 355902
rect 89798 355602 89824 355658
rect 90170 355602 90192 355658
rect 89798 355358 89824 355414
rect 90170 355358 90192 355414
rect 89798 355114 89824 355170
rect 90170 355114 90192 355170
rect 89798 354870 89824 354926
rect 90170 354870 90192 354926
rect 89798 354626 89824 354682
rect 90170 354626 90192 354682
rect 89798 354382 89824 354438
rect 90170 354382 90192 354438
rect 89798 354138 89824 354194
rect 90170 354138 90192 354194
rect 89798 353894 89824 353950
rect 90170 353894 90192 353950
rect 89432 149992 89488 150032
rect 89558 317350 89614 317390
rect 89558 149966 89614 317294
rect 89558 149870 89614 149910
rect 89810 317106 89866 317146
rect 89684 149844 89740 149884
rect 89684 147770 89740 149788
rect 89810 149722 89866 317050
rect 89810 149626 89866 149666
rect 89936 316862 89992 316902
rect 89936 149600 89992 316806
rect 90188 198684 90244 198724
rect 89936 149504 89992 149544
rect 90062 198440 90118 198480
rect 90062 149478 90118 198384
rect 90062 149382 90118 149422
rect 90188 149356 90244 198628
rect 90188 149260 90244 149300
rect 90314 198196 90370 198236
rect 90314 149234 90370 198140
rect 90314 149138 90370 149178
rect 89684 147704 89740 147714
rect 90468 147532 90524 365118
rect 93380 359562 93436 374257
rect 93380 359466 93436 359506
rect 110180 374927 110236 374976
rect 110180 359318 110236 374257
rect 110180 359222 110236 359262
rect 126980 374927 127036 374976
rect 126980 359074 127036 374257
rect 126980 358978 127036 359018
rect 143780 374927 143836 374976
rect 143780 358830 143836 374257
rect 200580 374927 200636 374976
rect 143780 358734 143836 358774
rect 199304 370786 199360 370826
rect 199304 357228 199360 370730
rect 200580 358586 200636 374257
rect 217380 374927 217436 374976
rect 200580 358490 200636 358530
rect 206864 370542 206920 370582
rect 206864 357228 206920 370486
rect 209258 370298 209314 370338
rect 209258 357228 209314 370242
rect 217380 358342 217436 374257
rect 244180 374927 244236 374976
rect 217380 358246 217436 358286
rect 229796 370054 229852 370094
rect 229796 357228 229852 369998
rect 230048 369810 230104 369850
rect 230048 357228 230104 369754
rect 232694 369566 232750 369606
rect 232694 357228 232750 369510
rect 232946 369322 233002 369362
rect 232946 357228 233002 369266
rect 233198 369078 233254 369118
rect 233198 357228 233254 369022
rect 241514 368834 241570 368874
rect 241514 357188 241570 368778
rect 244180 358098 244236 374257
rect 244180 358002 244236 358042
rect 260980 374927 261036 374976
rect 260980 357854 261036 374257
rect 277780 374927 277836 374976
rect 260980 357758 261036 357798
rect 266966 368590 267022 368630
rect 266966 357188 267022 368534
rect 268352 368346 268408 368386
rect 268100 365906 268156 365926
rect 268100 362001 268156 365850
rect 268100 361920 268156 361945
rect 268352 357188 268408 368290
rect 268604 368102 268660 368142
rect 268604 357188 268660 368046
rect 268856 367858 268912 367898
rect 268856 357188 268912 367802
rect 269108 367614 269164 367654
rect 269108 357188 269164 367558
rect 269360 367370 269416 367410
rect 269360 357188 269416 367314
rect 269612 367126 269668 367166
rect 269612 357188 269668 367070
rect 269864 366882 269920 366922
rect 269864 357188 269920 366826
rect 270116 366638 270172 366678
rect 270116 357188 270172 366582
rect 270368 366394 270424 366434
rect 270368 357188 270424 366338
rect 270620 366150 270676 366190
rect 270620 357188 270676 366094
rect 270872 365906 270928 365946
rect 270872 357188 270928 365850
rect 271124 365662 271180 365702
rect 271124 357188 271180 365606
rect 271376 365418 271432 365458
rect 271376 357188 271432 365362
rect 271628 365174 271684 365214
rect 271628 357188 271684 365118
rect 271880 364930 271936 364970
rect 271880 357188 271936 364874
rect 272132 364686 272188 364726
rect 272132 357188 272188 364630
rect 272384 364442 272440 364482
rect 272384 357188 272440 364386
rect 272636 364198 272692 364238
rect 272636 357648 272692 364142
rect 272636 357188 272692 357390
rect 272888 363954 272944 363994
rect 272888 357648 272944 363898
rect 272888 357188 272944 357390
rect 273140 363710 273196 363750
rect 273140 357648 273196 363654
rect 273140 357188 273196 357390
rect 273392 363466 273448 363506
rect 273392 357648 273448 363410
rect 273392 357188 273448 357390
rect 273644 363222 273700 363262
rect 273644 357648 273700 363166
rect 273644 357188 273700 357390
rect 273896 362978 273952 363018
rect 273896 357648 273952 362922
rect 273896 357188 273952 357390
rect 274148 362734 274204 362774
rect 274148 357648 274204 362678
rect 274148 357188 274204 357390
rect 274400 362490 274456 362530
rect 274400 357188 274456 362434
rect 274904 362490 274960 362530
rect 274652 362246 274708 362286
rect 274652 357188 274708 362190
rect 274904 357188 274960 362434
rect 275156 361758 275212 361798
rect 275156 357188 275212 361702
rect 275408 361514 275464 361554
rect 275408 357188 275464 361458
rect 277780 357610 277836 374257
rect 427200 374200 427400 375800
rect 441800 374200 442000 375800
rect 427200 374000 442000 374200
rect 444000 375800 458800 376000
rect 444000 374200 444200 375800
rect 458600 374200 458800 375800
rect 444000 374000 458800 374200
rect 466800 375800 481600 376000
rect 466800 374200 467000 375800
rect 481400 374200 481600 375800
rect 466800 374000 481600 374200
rect 470200 373500 470900 373600
rect 470200 373000 470300 373500
rect 470800 373000 470900 373500
rect 470200 372900 470900 373000
rect 471400 373500 472100 373600
rect 471400 373000 471500 373500
rect 472000 373000 472100 373500
rect 471400 372900 472100 373000
rect 480662 370636 480718 370676
rect 320670 365486 322812 365612
rect 320670 364604 320796 365486
rect 322686 364604 322812 365486
rect 328500 365400 329300 365500
rect 328500 364800 328600 365400
rect 329200 364800 329300 365400
rect 328500 364700 329300 364800
rect 320670 364478 322812 364604
rect 328500 364000 329300 364100
rect 319645 363600 319701 363621
rect 277780 357514 277836 357554
rect 292040 362734 292096 362774
rect 292040 357188 292096 362678
rect 292292 362490 292348 362530
rect 292292 357188 292348 362434
rect 309302 362246 309358 362286
rect 309302 357188 309358 362190
rect 309554 362002 309610 362042
rect 309554 357188 309610 361946
rect 309806 361758 309862 361798
rect 309806 357188 309862 361702
rect 310058 361514 310114 361554
rect 310058 357188 310114 361458
rect 319645 361422 319701 363544
rect 320684 363376 320740 363402
rect 320684 363034 320740 363320
rect 328500 363400 328600 364000
rect 329200 363400 329300 364000
rect 328500 363300 329300 363400
rect 472400 363600 478000 363800
rect 320996 362908 321020 362964
rect 321188 362908 321209 362964
rect 320684 362815 320740 362847
rect 321022 362244 321079 362908
rect 310310 361270 310366 361310
rect 319645 361238 319701 361252
rect 320668 362184 321079 362244
rect 321930 362502 323442 362628
rect 310310 357188 310366 361214
rect 310562 361026 310618 361066
rect 310562 357188 310618 360970
rect 316764 360990 317772 361116
rect 310814 360782 310870 360822
rect 310814 357188 310870 360726
rect 316764 360612 316890 360990
rect 317646 360612 317772 360990
rect 311066 360538 311122 360578
rect 316764 360486 317772 360612
rect 311066 357188 311122 360482
rect 311318 360294 311374 360334
rect 311318 357188 311374 360238
rect 311570 360050 311626 360090
rect 311570 357188 311626 359994
rect 311822 359806 311878 359846
rect 311822 357188 311878 359750
rect 312074 359562 312130 359778
rect 312074 357188 312130 359506
rect 312326 359318 312382 359778
rect 312326 357188 312382 359262
rect 312578 359074 312634 359778
rect 312578 357188 312634 359018
rect 312830 358830 312886 359778
rect 312830 357188 312886 358774
rect 313082 358586 313138 359778
rect 313082 357188 313138 358530
rect 313334 358342 313390 359778
rect 313334 357188 313390 358286
rect 313586 358098 313642 359778
rect 313586 357188 313642 358042
rect 313838 357854 313894 359778
rect 313838 357188 313894 357798
rect 314090 357610 314146 359778
rect 314090 357188 314146 357554
rect 314342 359074 314398 359778
rect 314342 357188 314398 359018
rect 314594 358830 314650 359778
rect 314594 357188 314650 358774
rect 314846 358586 314902 359778
rect 314846 357188 314902 358530
rect 315098 358342 315154 359778
rect 315098 357188 315154 358286
rect 315350 358098 315406 359778
rect 315350 357188 315406 358042
rect 315602 357854 315658 359778
rect 315602 357188 315658 357798
rect 315854 357610 315910 359778
rect 320668 359647 320728 362184
rect 321930 361872 322056 362502
rect 323316 361872 323442 362502
rect 321930 361746 323442 361872
rect 334400 362200 346200 362400
rect 321040 361525 321096 361565
rect 321040 360559 321096 361265
rect 334400 360800 334600 362200
rect 346000 360800 346200 362200
rect 334400 360600 346200 360800
rect 320908 360499 321096 360559
rect 320908 359647 320968 360499
rect 315854 357188 315910 357554
rect 472400 349200 472600 363600
rect 477800 349200 478000 363600
rect 472400 349000 478000 349200
rect 410640 342436 410700 342904
rect 410640 342340 410700 342380
rect 410800 342310 410860 342904
rect 410800 342216 410860 342254
rect 410130 341712 412020 341838
rect 410130 340578 410256 341712
rect 411894 340578 412020 341712
rect 410130 340452 412020 340578
rect 396116 339676 396172 339696
rect 389438 332356 389494 332396
rect 385658 332112 385714 332152
rect 381878 331868 381934 331908
rect 378098 331624 378154 331664
rect 374318 331380 374374 331420
rect 370538 331136 370594 331176
rect 366758 330892 366814 330932
rect 363104 330648 363160 330688
rect 359324 330404 359380 330444
rect 355544 330160 355600 330200
rect 351764 329916 351820 329956
rect 347984 329672 348040 329712
rect 344204 329428 344260 329468
rect 340424 329184 340480 329224
rect 336644 328940 336700 328980
rect 332990 328696 333046 328736
rect 332990 316862 333046 328640
rect 316358 316798 316414 316834
rect 332990 316655 333046 316684
rect 333368 327720 333424 327760
rect 333368 316862 333424 327664
rect 333368 316655 333424 316684
rect 333872 324548 333928 324588
rect 333872 316862 333928 324492
rect 333872 316655 333928 316684
rect 336644 316862 336700 328884
rect 336644 316655 336700 316684
rect 337148 327720 337204 327760
rect 337148 316862 337204 327664
rect 337148 316655 337204 316684
rect 337652 324304 337708 324344
rect 337652 316862 337708 324248
rect 337652 316655 337708 316684
rect 340424 316862 340480 329128
rect 340424 316655 340480 316684
rect 340928 327720 340984 327760
rect 340928 316862 340984 327664
rect 340928 316655 340984 316684
rect 341432 324060 341488 324100
rect 341432 316862 341488 324004
rect 341432 316655 341488 316684
rect 344204 316862 344260 329372
rect 344204 316655 344260 316684
rect 344708 327720 344764 327760
rect 344708 316862 344764 327664
rect 344708 316655 344764 316684
rect 345212 323816 345268 323856
rect 345212 316862 345268 323760
rect 345212 316655 345268 316684
rect 347984 316862 348040 329616
rect 347984 316655 348040 316684
rect 348488 327720 348544 327760
rect 348488 316862 348544 327664
rect 348488 316655 348544 316684
rect 348992 323572 349048 323612
rect 348992 316862 349048 323516
rect 348992 316655 349048 316684
rect 351764 316862 351820 329860
rect 351764 316655 351820 316684
rect 352268 327720 352324 327760
rect 352268 316862 352324 327664
rect 352268 316655 352324 316684
rect 352772 323328 352828 323368
rect 352772 316862 352828 323272
rect 352772 316655 352828 316684
rect 355544 316862 355600 330104
rect 355544 316655 355600 316684
rect 356048 327720 356104 327760
rect 356048 316862 356104 327664
rect 356048 316655 356104 316684
rect 356552 323084 356608 323124
rect 356552 316862 356608 323028
rect 356552 316655 356608 316684
rect 359324 316862 359380 330348
rect 359324 316655 359380 316684
rect 359828 327720 359884 327760
rect 359828 316862 359884 327664
rect 359828 316655 359884 316684
rect 360332 322840 360388 322880
rect 360332 316862 360388 322784
rect 360332 316655 360388 316684
rect 363104 316862 363160 330592
rect 363104 316655 363160 316684
rect 363608 327964 363664 328004
rect 363608 316862 363664 327908
rect 363608 316655 363664 316684
rect 364112 322596 364168 322636
rect 364112 316862 364168 322540
rect 364112 316655 364168 316684
rect 366758 316862 366814 330836
rect 366758 316655 366814 316684
rect 367262 327964 367318 328004
rect 367262 316862 367318 327908
rect 367262 316655 367318 316684
rect 367766 322352 367822 322392
rect 367766 316862 367822 322296
rect 367766 316655 367822 316684
rect 370538 316862 370594 331080
rect 370538 316655 370594 316684
rect 371042 327964 371098 328004
rect 371042 316862 371098 327908
rect 371042 316655 371098 316684
rect 371546 322108 371602 322148
rect 371546 316862 371602 322052
rect 371546 316655 371602 316684
rect 374318 316862 374374 331324
rect 374318 316655 374374 316684
rect 374822 327964 374878 328004
rect 374822 316862 374878 327908
rect 374822 316655 374878 316684
rect 375326 321864 375382 321904
rect 375326 316862 375382 321808
rect 375326 316655 375382 316684
rect 378098 316862 378154 331568
rect 378098 316655 378154 316684
rect 378602 327964 378658 328004
rect 378602 316862 378658 327908
rect 378602 316655 378658 316684
rect 379106 321620 379162 321660
rect 379106 316862 379162 321564
rect 379106 316655 379162 316684
rect 381878 316862 381934 331812
rect 381878 316655 381934 316684
rect 382382 327964 382438 328004
rect 382382 316862 382438 327908
rect 382382 316655 382438 316684
rect 382886 321376 382942 321416
rect 382886 316862 382942 321320
rect 382886 316655 382942 316684
rect 385658 316862 385714 332056
rect 385658 316655 385714 316684
rect 386162 327964 386218 328004
rect 386162 316862 386218 327908
rect 386162 316655 386218 316684
rect 386666 321132 386722 321172
rect 386666 316862 386722 321076
rect 386666 316655 386722 316684
rect 389438 316862 389494 332300
rect 389438 316655 389494 316684
rect 389942 327964 389998 328004
rect 389942 316862 389998 327908
rect 389942 316655 389998 316684
rect 390446 320888 390502 320928
rect 390446 316862 390502 320832
rect 395612 316862 395668 316902
rect 396116 316862 396172 339620
rect 465290 336260 465346 336300
rect 461510 336016 461566 336056
rect 457730 335772 457786 335812
rect 454076 335528 454132 335568
rect 450296 335284 450352 335324
rect 446516 335040 446572 335080
rect 442736 334796 442792 334836
rect 438956 334552 439012 334592
rect 435176 334308 435232 334348
rect 431396 334064 431452 334104
rect 427616 333820 427672 333860
rect 423962 333576 424018 333616
rect 420182 333332 420238 333372
rect 416402 333088 416458 333128
rect 412622 332844 412678 332884
rect 408842 332600 408898 332640
rect 404558 327476 404614 327516
rect 404054 327232 404110 327272
rect 401534 326988 401590 327028
rect 395540 316684 395558 316740
rect 395714 316684 395732 316740
rect 390446 316655 390502 316684
rect 395612 316655 395668 316684
rect 396116 316655 396172 316684
rect 396872 326744 396928 326784
rect 396872 316862 396928 326688
rect 396872 316655 396928 316684
rect 398006 326500 398062 326540
rect 398006 316862 398062 326444
rect 398006 316655 398062 316684
rect 401534 316862 401590 326932
rect 402542 326256 402598 326296
rect 401534 316655 401590 316684
rect 402038 326012 402094 326052
rect 402038 316862 402094 325956
rect 402038 316655 402094 316684
rect 402542 316862 402598 326200
rect 402542 316655 402598 316684
rect 403046 325768 403102 325808
rect 403046 316862 403102 325712
rect 403046 316655 403102 316684
rect 403550 325524 403606 325564
rect 403550 316862 403606 325468
rect 403550 316655 403606 316684
rect 404054 316862 404110 327176
rect 404054 316655 404110 316684
rect 404558 316862 404614 327420
rect 404558 316655 404614 316684
rect 405062 325280 405118 325320
rect 405062 316862 405118 325224
rect 405062 316655 405118 316684
rect 405566 325036 405622 325076
rect 405566 316862 405622 324980
rect 405566 316655 405622 316684
rect 406070 324792 406126 324832
rect 406070 316862 406126 324736
rect 406070 316655 406126 316684
rect 408842 316862 408898 332544
rect 408842 316655 408898 316684
rect 409346 328208 409402 328248
rect 409346 316862 409402 328152
rect 409346 316655 409402 316684
rect 409850 320644 409906 320684
rect 409850 316862 409906 320588
rect 409850 316655 409906 316684
rect 412622 316862 412678 332788
rect 412622 316655 412678 316684
rect 413126 328208 413182 328248
rect 413126 316862 413182 328152
rect 413126 316655 413182 316684
rect 413630 320400 413686 320440
rect 413630 316862 413686 320344
rect 413630 316655 413686 316684
rect 416402 316862 416458 333032
rect 416402 316655 416458 316684
rect 416906 328208 416962 328248
rect 416906 316862 416962 328152
rect 416906 316655 416962 316684
rect 417410 320156 417466 320196
rect 417410 316862 417466 320100
rect 417410 316655 417466 316684
rect 420182 316862 420238 333276
rect 420182 316655 420238 316684
rect 420686 328208 420742 328248
rect 420686 316862 420742 328152
rect 420686 316655 420742 316684
rect 421190 319912 421246 319952
rect 421190 316862 421246 319856
rect 421190 316655 421246 316684
rect 423962 316862 424018 333520
rect 423962 316655 424018 316684
rect 424466 328208 424522 328248
rect 424466 316862 424522 328152
rect 424466 316655 424522 316684
rect 424970 319668 425026 319708
rect 424970 316862 425026 319612
rect 424970 316655 425026 316684
rect 427616 316862 427672 333764
rect 427616 316655 427672 316684
rect 428120 328208 428176 328248
rect 428120 316862 428176 328152
rect 428120 316655 428176 316684
rect 428624 319424 428680 319464
rect 428624 316862 428680 319368
rect 428624 316655 428680 316684
rect 431396 316862 431452 334008
rect 431396 316655 431452 316684
rect 431900 328208 431956 328248
rect 431900 316862 431956 328152
rect 431900 316655 431956 316684
rect 432404 319180 432460 319220
rect 432404 316862 432460 319124
rect 432404 316655 432460 316684
rect 435176 316862 435232 334252
rect 435176 316655 435232 316684
rect 435680 328208 435736 328248
rect 435680 316862 435736 328152
rect 435680 316655 435736 316684
rect 436184 318936 436240 318976
rect 436184 316862 436240 318880
rect 436184 316655 436240 316684
rect 438956 316862 439012 334496
rect 438956 316655 439012 316684
rect 439460 328452 439516 328492
rect 439460 316862 439516 328396
rect 439460 316655 439516 316684
rect 439964 318692 440020 318732
rect 439964 316862 440020 318636
rect 439964 316655 440020 316684
rect 442736 316862 442792 334740
rect 442736 316655 442792 316684
rect 443240 328452 443296 328492
rect 443240 316862 443296 328396
rect 443240 316655 443296 316684
rect 443744 318448 443800 318488
rect 443744 316862 443800 318392
rect 443744 316655 443800 316684
rect 446516 316862 446572 334984
rect 446516 316655 446572 316684
rect 447020 328452 447076 328492
rect 447020 316862 447076 328396
rect 447020 316655 447076 316684
rect 447524 318204 447580 318244
rect 447524 316862 447580 318148
rect 447524 316655 447580 316684
rect 450296 316862 450352 335228
rect 450296 316655 450352 316684
rect 450800 328452 450856 328492
rect 450800 316862 450856 328396
rect 450800 316655 450856 316684
rect 451304 317960 451360 318000
rect 451304 316862 451360 317904
rect 451304 316655 451360 316684
rect 454076 316862 454132 335472
rect 454076 316655 454132 316684
rect 454580 328452 454636 328492
rect 454580 316862 454636 328396
rect 454580 316655 454636 316684
rect 455084 317716 455140 317756
rect 455084 316862 455140 317660
rect 455084 316655 455140 316684
rect 457730 316862 457786 335716
rect 457730 316655 457786 316684
rect 458234 328452 458290 328492
rect 458234 316862 458290 328396
rect 458234 316655 458290 316684
rect 458738 317472 458794 317512
rect 458738 316862 458794 317416
rect 458738 316655 458794 316684
rect 461510 316862 461566 335960
rect 461510 316655 461566 316684
rect 462014 328452 462070 328492
rect 462014 316862 462070 328396
rect 462014 316655 462070 316684
rect 462518 317228 462574 317268
rect 462518 316862 462574 317172
rect 462518 316655 462574 316684
rect 465290 316862 465346 336204
rect 477548 332524 477644 332542
rect 477548 332192 477644 332418
rect 477548 332054 477644 332080
rect 477862 332528 477984 349000
rect 480410 339508 480466 339548
rect 480158 339264 480214 339304
rect 479906 339020 479962 339060
rect 479654 338776 479710 338816
rect 479402 338532 479458 338572
rect 479150 338288 479206 338328
rect 478898 338004 478954 338044
rect 477552 331596 477648 331632
rect 477552 331092 477648 331474
rect 477552 330970 477648 330986
rect 477862 331104 477984 332400
rect 465290 316655 465346 316684
rect 465794 328452 465850 328492
rect 465794 316862 465850 328396
rect 465794 316655 465850 316684
rect 466298 316984 466354 317024
rect 466298 316862 466354 316928
rect 466298 316655 466354 316684
rect 201194 147648 201250 148624
rect 90468 147466 90524 147476
rect 115668 147532 115724 147542
rect 88424 147334 88480 147364
rect 88046 146626 88480 146682
rect 86968 137700 87024 137710
rect 86282 130551 86338 130577
rect 88424 109928 88480 146626
rect 89152 139328 90832 139440
rect 89152 138432 89264 139328
rect 90720 138432 90832 139328
rect 89152 138320 90832 138432
rect 115668 139244 115724 147476
rect 126644 147526 126700 147566
rect 117012 147308 117068 147335
rect 116787 147084 116843 147104
rect 115220 123452 115276 123462
rect 90342 110880 90972 111006
rect 90342 110502 90468 110880
rect 90846 110502 90972 110880
rect 115220 110908 115276 123396
rect 115387 123217 115443 123231
rect 115387 111126 115443 123161
rect 115668 111388 115725 139244
rect 115892 138254 115948 138294
rect 115892 111612 115948 138198
rect 116116 138132 116172 138172
rect 116116 111836 116172 138076
rect 116564 138010 116620 138050
rect 116340 137888 116396 137928
rect 116340 113068 116396 137832
rect 116564 114076 116620 137954
rect 116564 113980 116620 114020
rect 116340 112928 116396 113012
rect 116116 111780 116620 111836
rect 115892 111556 116396 111612
rect 115668 111332 116173 111388
rect 115387 111070 115905 111126
rect 115220 110852 115724 110908
rect 90342 110376 90972 110502
rect 88424 109858 89510 109928
rect 86412 109620 86640 109646
rect 86412 108738 86640 109368
rect 86412 108524 86640 108538
rect 80836 108486 80892 108500
rect 86650 108162 86950 108238
rect 74214 107856 75222 107982
rect 74214 107352 74340 107856
rect 75096 107352 75222 107856
rect 74214 107226 75222 107352
rect 86650 107072 86726 108162
rect 90342 107982 90594 110376
rect 91350 109620 91854 109746
rect 91350 108738 91476 109620
rect 91728 108738 91854 109620
rect 91350 108612 91854 108738
rect 90342 107856 90972 107982
rect 90342 107478 90468 107856
rect 90846 107478 90972 107856
rect 90342 107352 90972 107478
rect 92358 107856 93114 107982
rect 92358 107352 92484 107856
rect 92988 107352 93114 107856
rect 92358 107226 93114 107352
rect 74050 107016 74074 107072
rect 74196 107016 86726 107072
rect 73472 106676 73528 106690
rect 77864 106907 77932 106925
rect 68436 106198 68450 106254
rect 68678 106198 68692 106254
rect 71652 106228 71708 106248
rect 77696 106304 77764 106344
rect 77696 105957 77764 106248
rect 77864 105957 77932 106755
rect 102081 106907 102141 106927
rect 102081 106068 102141 106755
rect 102481 106907 102541 106921
rect 102281 106605 102341 106623
rect 102281 106068 102341 106453
rect 102481 106068 102541 106755
rect 102681 106605 102741 106627
rect 102681 106068 102741 106453
rect 103068 106452 103100 106508
rect 103156 106452 107641 106508
rect 107581 106050 107641 106452
rect 102081 83802 102141 84121
rect 102281 83802 102341 84121
rect 102481 83802 102541 84121
rect 102681 83802 102741 84121
rect 107581 83906 107641 84118
rect 35524 78054 35580 78102
rect 115668 78012 115724 110852
rect 32550 75674 32606 75734
rect 32550 32680 32606 75374
rect 32802 75674 32858 75734
rect 32802 33176 32858 75374
rect 33054 75674 33110 75734
rect 33054 33428 33110 75374
rect 33306 75674 33362 75734
rect 33306 33680 33362 75374
rect 33558 75674 33614 75734
rect 33558 33932 33614 75374
rect 33810 75674 33866 75734
rect 33810 34184 33866 75374
rect 115668 75404 115724 77956
rect 115668 75338 115724 75348
rect 115849 74749 115905 111070
rect 115849 74683 115905 74693
rect 114597 72198 115227 72261
rect 113148 72072 114030 72198
rect 112494 71868 112570 71906
rect 112494 70113 112570 71588
rect 113148 71442 113274 72072
rect 113904 71442 114030 72072
rect 114597 71694 114660 72198
rect 115164 71694 115227 72198
rect 114597 71631 115227 71694
rect 116117 71620 116173 111332
rect 116340 81932 116396 111556
rect 116340 81836 116396 81876
rect 116564 80700 116620 111780
rect 116564 80604 116620 80644
rect 116787 72660 116843 147028
rect 117012 72820 117068 147252
rect 117460 143622 117516 143668
rect 117236 138376 117292 138398
rect 117236 112060 117292 138320
rect 117460 126844 117516 143566
rect 117460 126748 117516 126788
rect 117684 143500 117740 143540
rect 117684 125836 117740 143444
rect 117684 125740 117740 125780
rect 117908 143378 117964 143418
rect 117908 119900 117964 143322
rect 117908 119804 117964 119844
rect 118132 143256 118188 143296
rect 118132 119004 118188 143200
rect 118132 118908 118188 118948
rect 118356 143134 118412 143174
rect 118132 118668 118188 118708
rect 117908 118444 117964 118484
rect 117684 118220 117740 118260
rect 117236 111956 117292 112004
rect 117460 117996 117516 118036
rect 117460 111500 117516 117940
rect 117460 111404 117516 111444
rect 117684 110044 117740 118164
rect 117684 109948 117740 109988
rect 117908 108504 117964 118388
rect 117908 108408 117964 108448
rect 118132 107048 118188 118612
rect 118356 117996 118412 143078
rect 118356 117900 118412 117940
rect 118580 143012 118636 143052
rect 118580 116988 118636 142956
rect 118580 116892 118636 116932
rect 118804 142890 118860 142930
rect 118804 115980 118860 142834
rect 118804 115884 118860 115924
rect 119028 142768 119084 142808
rect 119028 114972 119084 142712
rect 125524 138742 125580 138782
rect 123620 138620 123676 138660
rect 123620 128574 123676 138564
rect 124628 137368 124684 137387
rect 124628 128574 124684 137312
rect 125524 128574 125580 138686
rect 125860 138498 125916 138538
rect 125860 128574 125916 138442
rect 126644 128574 126700 147470
rect 128884 147404 128940 147444
rect 126980 142646 127036 142686
rect 126980 128574 127036 142590
rect 128884 128574 128940 147348
rect 131124 147282 131180 147322
rect 201194 147254 201250 147592
rect 129220 142524 129276 142564
rect 129220 128574 129276 142468
rect 131124 128574 131180 147226
rect 133364 147160 133420 147200
rect 131460 142402 131516 142442
rect 131460 128574 131516 142346
rect 133364 128574 133420 147104
rect 135604 147038 135660 147078
rect 133700 142280 133756 142320
rect 133700 128574 133756 142224
rect 135604 128574 135660 146982
rect 137844 146916 137900 146956
rect 135940 142158 135996 142198
rect 135940 128574 135996 142102
rect 137844 128574 137900 146860
rect 140084 146794 140140 146834
rect 138180 142036 138236 142076
rect 138180 128574 138236 141980
rect 140084 128574 140140 146738
rect 142324 146672 142380 146712
rect 140420 141914 140476 141954
rect 140420 128574 140476 141858
rect 142324 128574 142380 146616
rect 145012 146550 145068 146590
rect 142660 141792 142716 141832
rect 142660 128574 142716 141736
rect 145012 128574 145068 146494
rect 147252 146428 147308 146468
rect 145348 141670 145404 141710
rect 145348 128574 145404 141614
rect 147252 128574 147308 146372
rect 149492 146306 149548 146346
rect 147588 141548 147644 141588
rect 147588 128574 147644 141492
rect 149492 128574 149548 146250
rect 151732 146184 151788 146224
rect 149828 141426 149884 141466
rect 149828 128574 149884 141370
rect 151732 128574 151788 146128
rect 153972 146062 154028 146102
rect 152068 141304 152124 141344
rect 152068 128574 152124 141248
rect 153972 128574 154028 146006
rect 156212 145940 156268 145980
rect 154308 141182 154364 141222
rect 154308 128574 154364 141126
rect 156212 128574 156268 145884
rect 158452 145818 158508 145858
rect 156548 141060 156604 141100
rect 156548 128574 156604 141004
rect 158452 128574 158508 145762
rect 160692 145696 160748 145736
rect 158788 140938 158844 140978
rect 158788 128574 158844 140882
rect 160692 128574 160748 145640
rect 163380 145574 163436 145614
rect 161028 140816 161084 140856
rect 161028 128574 161084 140760
rect 163380 128574 163436 145518
rect 165620 145452 165676 145492
rect 163716 140694 163772 140734
rect 163716 128574 163772 140638
rect 165620 128574 165676 145396
rect 167860 145330 167916 145370
rect 165956 140572 166012 140612
rect 165956 128574 166012 140516
rect 167860 128574 167916 145274
rect 170100 145208 170156 145248
rect 168196 140450 168252 140490
rect 168196 128574 168252 140394
rect 170100 128574 170156 145152
rect 172340 145086 172396 145126
rect 170436 140328 170492 140368
rect 170436 128574 170492 140272
rect 172340 128574 172396 145030
rect 174580 144964 174636 145004
rect 172676 140206 172732 140246
rect 172676 128574 172732 140150
rect 174580 128574 174636 144908
rect 176820 144842 176876 144882
rect 174916 140084 174972 140124
rect 174916 128574 174972 140028
rect 176820 128574 176876 144786
rect 179060 144720 179116 144760
rect 177156 139962 177212 140002
rect 177156 128574 177212 139906
rect 179060 128574 179116 144664
rect 181748 144598 181804 144638
rect 179396 139840 179452 139880
rect 179396 128574 179452 139784
rect 181748 128574 181804 144542
rect 183988 144476 184044 144516
rect 182084 139718 182140 139758
rect 182084 128574 182140 139662
rect 183988 128574 184044 144420
rect 186228 144354 186284 144394
rect 184324 139596 184380 139636
rect 184324 128574 184380 139540
rect 186228 128574 186284 144298
rect 188468 144232 188524 144272
rect 186564 139474 186620 139514
rect 186564 128574 186620 139418
rect 188468 128574 188524 144176
rect 190708 144110 190764 144150
rect 188804 139352 188860 139392
rect 188804 128574 188860 139296
rect 190708 128574 190764 144054
rect 192948 143988 193004 144028
rect 191044 139230 191100 139270
rect 191044 128574 191100 139174
rect 192948 128574 193004 143932
rect 195188 143866 195244 143906
rect 193284 139108 193340 139148
rect 193284 128574 193340 139052
rect 195188 128574 195244 143810
rect 197428 143744 197484 143784
rect 195524 138986 195580 139026
rect 195524 128574 195580 138930
rect 197428 128608 197484 143688
rect 197764 138864 197820 138904
rect 197764 128608 197820 138808
rect 202328 129379 202384 148624
rect 202580 147892 202636 148624
rect 202580 147254 202636 147836
rect 202832 148136 202888 148624
rect 202832 147254 202888 148080
rect 202328 129041 202384 129086
rect 203084 129380 203140 148624
rect 203084 129041 203140 129075
rect 203336 129385 203392 148624
rect 203336 129041 203392 129062
rect 203588 129372 203644 148624
rect 203588 129041 203644 129064
rect 203840 129370 203896 148624
rect 214172 148258 214228 148625
rect 214172 148162 214228 148202
rect 233610 148014 233666 148665
rect 233610 147864 233666 147958
rect 292670 148258 292726 148268
rect 203840 129041 203896 129061
rect 206990 137368 207046 137378
rect 201663 120593 205130 120831
rect 204892 118890 205130 120593
rect 206990 120204 207046 137312
rect 275800 133700 276600 133800
rect 275800 133100 275900 133700
rect 276500 133100 276600 133700
rect 275800 133000 276600 133100
rect 275800 132300 276600 132400
rect 275800 131700 275900 132300
rect 276500 131700 276600 132300
rect 275800 131600 276600 131700
rect 206990 119672 207046 119700
rect 204892 118652 207888 118890
rect 119028 114876 119084 114916
rect 118132 106952 118188 106992
rect 201658 87317 207858 87551
rect 201662 86516 207866 86598
rect 201639 86316 207898 86398
rect 201639 86116 207898 86198
rect 201639 85916 207898 85998
rect 201639 85716 207898 85798
rect 201639 85506 207898 85588
rect 201639 85296 207898 85378
rect 201639 85086 207898 85168
rect 201639 84876 207898 84958
rect 201639 84674 207898 84756
rect 201639 84476 207898 84558
rect 201639 84270 207898 84352
rect 201639 84066 207898 84148
rect 201639 83862 207898 83944
rect 201639 83658 207898 83740
rect 201639 83454 207898 83536
rect 201639 83250 207898 83332
rect 201639 83046 207898 83128
rect 201658 80551 207873 80630
rect 201639 80347 207898 80426
rect 201639 80143 207898 80222
rect 201639 79883 207898 79962
rect 201656 78805 207866 79336
rect 206990 78624 207046 78652
rect 202328 78411 202384 78439
rect 122052 75488 122108 75804
rect 122388 75404 122444 75804
rect 122388 75338 122444 75348
rect 124404 75404 124460 75804
rect 124404 75338 124460 75348
rect 126420 74749 126476 75804
rect 128436 75404 128492 75804
rect 128436 75338 128492 75348
rect 126420 74683 126476 74693
rect 135946 72828 140986 72954
rect 117012 72760 119264 72820
rect 119904 72760 134560 72820
rect 116787 72600 119264 72660
rect 119904 72600 134400 72660
rect 117465 71802 117541 71824
rect 116038 71564 116067 71620
rect 116239 71564 116272 71620
rect 117465 71614 117470 71802
rect 117534 71614 117541 71802
rect 113148 71316 114030 71442
rect 117465 70844 117541 71614
rect 117465 70768 129798 70844
rect 117465 70766 117541 70768
rect 129722 70126 129798 70768
rect 134340 70680 134400 72600
rect 134500 70680 134560 72760
rect 135946 71442 136072 72828
rect 140860 71442 140986 72828
rect 135946 71316 140986 71442
rect 34400 57600 36400 57800
rect 34400 43200 34600 57600
rect 36200 43200 36400 57600
rect 202328 54452 202384 78126
rect 203084 78404 203140 78439
rect 203084 54720 203140 78128
rect 203336 78404 203392 78439
rect 203336 54972 203392 78128
rect 203588 78404 203644 78439
rect 203588 55224 203644 78128
rect 203840 78404 203896 78439
rect 203840 55476 203896 78128
rect 206990 61768 207046 78120
rect 207579 75348 207589 75404
rect 207645 75348 207655 75404
rect 207589 62081 207645 75348
rect 207589 62025 218290 62081
rect 206990 61712 208656 61768
rect 208801 61712 208826 61768
rect 204957 59840 213764 59885
rect 204957 59033 205006 59840
rect 206669 59033 213764 59840
rect 204957 58998 213764 59033
rect 213886 58998 213966 59885
rect 203840 55420 217576 55476
rect 203588 55168 217324 55224
rect 203336 54916 217072 54972
rect 203084 54664 216820 54720
rect 202328 54396 216568 54452
rect 199000 53800 204646 54000
rect 199000 51600 199200 53800
rect 204464 51600 204646 53800
rect 199000 51400 204646 51600
rect 205266 53800 211000 54000
rect 205266 51600 205440 53800
rect 210800 51600 211000 53800
rect 205266 51400 211000 51600
rect 34400 43000 36400 43200
rect 59700 41700 60500 41800
rect 59700 41100 59800 41700
rect 60400 41100 60500 41700
rect 59700 41000 60500 41100
rect 59700 40500 60500 40600
rect 59700 39900 59800 40500
rect 60400 39900 60500 40500
rect 59700 39800 60500 39900
rect 102200 35400 117000 35600
rect 33810 34128 34992 34184
rect 35048 34128 35088 34184
rect 33558 33876 34362 33932
rect 34418 33876 34458 33932
rect 102200 33800 102400 35400
rect 116800 33800 117000 35400
rect 33306 33624 73422 33680
rect 73478 33624 73518 33680
rect 102200 33600 117000 33800
rect 216512 33662 216568 54396
rect 216764 33930 216820 54664
rect 217016 34182 217072 54916
rect 217268 34434 217324 55168
rect 217520 34686 217576 55420
rect 218234 34969 218290 62025
rect 292670 61630 292726 148202
rect 292922 148014 292978 148054
rect 292922 61882 292978 147958
rect 293174 62134 293230 148624
rect 293426 62386 293482 148596
rect 293678 62638 293734 148596
rect 293930 62890 293986 148596
rect 294182 63142 294238 148596
rect 294434 63394 294490 148596
rect 294686 63646 294742 148596
rect 294938 63898 294994 148596
rect 295190 64150 295246 148596
rect 295442 64402 295498 148596
rect 295694 147770 295750 148596
rect 295694 146644 295750 147714
rect 295946 137888 296002 148596
rect 296198 138010 296254 148596
rect 296450 138132 296506 148596
rect 296702 138254 296758 148596
rect 296954 138376 297010 148596
rect 297206 138498 297262 148596
rect 297458 138620 297514 148596
rect 297710 138742 297766 148596
rect 297962 138864 298018 148596
rect 298214 138986 298270 148596
rect 298466 139108 298522 148596
rect 298718 139230 298774 148596
rect 298970 139352 299026 148596
rect 299222 139474 299278 148596
rect 299474 139596 299530 148596
rect 299726 139718 299782 148596
rect 299978 139840 300034 148596
rect 300230 139962 300286 148596
rect 300482 140084 300538 148596
rect 300734 140206 300790 148596
rect 300986 140328 301042 148596
rect 301238 140450 301294 148596
rect 301490 140572 301546 148596
rect 301742 140694 301798 148596
rect 301994 140816 302050 148596
rect 302246 140938 302302 148596
rect 302498 141060 302554 148596
rect 302750 141182 302806 148596
rect 303002 141304 303058 148596
rect 303254 141426 303310 148596
rect 303506 141548 303562 148596
rect 303758 141670 303814 148596
rect 304010 141792 304066 148596
rect 304262 141914 304318 148596
rect 304514 142036 304570 148596
rect 304766 142158 304822 148596
rect 305018 142280 305074 148596
rect 305270 142402 305326 148596
rect 305522 142524 305578 148596
rect 305774 142646 305830 148596
rect 306026 142768 306082 148596
rect 306278 142890 306334 148596
rect 306530 143012 306586 148596
rect 306782 143134 306838 148596
rect 307034 143256 307090 148596
rect 307286 143378 307342 148596
rect 307538 143500 307594 148596
rect 307790 143622 307846 148596
rect 308042 143744 308098 148596
rect 308294 143866 308350 148596
rect 308546 143988 308602 148596
rect 308798 144110 308854 148596
rect 309050 144232 309106 148596
rect 309302 144354 309358 148596
rect 309554 144476 309610 148596
rect 309806 144598 309862 148596
rect 310058 144720 310114 148596
rect 310310 144842 310366 148596
rect 310562 144964 310618 148596
rect 310814 145086 310870 148596
rect 311066 145208 311122 148596
rect 311318 145330 311374 148596
rect 311570 145452 311626 148596
rect 311822 145574 311878 148596
rect 312074 145696 312130 148596
rect 312326 145818 312382 148596
rect 312578 145940 312634 148596
rect 312830 146062 312886 148596
rect 313082 146184 313138 148596
rect 313334 146306 313390 148596
rect 313586 146428 313642 148596
rect 313838 146550 313894 148596
rect 314090 146672 314146 148596
rect 314342 146794 314398 148596
rect 314342 146698 314398 146738
rect 314594 146916 314650 148596
rect 314594 146701 314650 146860
rect 314846 147038 314902 148596
rect 314846 146701 314902 146982
rect 315098 147160 315154 148596
rect 315098 146701 315154 147104
rect 315350 147282 315406 148596
rect 315350 146701 315406 147226
rect 315602 147404 315658 148596
rect 315602 146701 315658 147348
rect 315854 147526 315910 148596
rect 316358 147892 316414 316615
rect 477548 315724 477644 315742
rect 477548 315392 477644 315618
rect 477548 315254 477644 315280
rect 477862 315728 477984 330976
rect 477552 314796 477648 314832
rect 477552 314292 477648 314674
rect 477552 314170 477648 314186
rect 477862 314304 477984 315600
rect 477548 298924 477644 298942
rect 477548 298592 477644 298818
rect 477548 298454 477644 298480
rect 477862 298928 477984 314176
rect 477552 297996 477648 298032
rect 477552 297492 477648 297874
rect 477552 297370 477648 297386
rect 477862 297504 477984 298800
rect 477548 225324 477644 225342
rect 477548 224992 477644 225218
rect 477548 224854 477644 224880
rect 477862 225328 477984 297376
rect 477552 224396 477648 224432
rect 477552 223892 477648 224274
rect 477552 223770 477648 223786
rect 477862 223904 477984 225200
rect 478646 337760 478702 337800
rect 478646 224358 478702 337704
rect 478898 246562 478954 337948
rect 478898 246400 478954 246440
rect 478646 224196 478702 224236
rect 477862 223359 477984 223776
rect 321000 149736 321600 149836
rect 321000 149336 321100 149736
rect 321500 149336 321600 149736
rect 321000 149236 321600 149336
rect 321000 148736 321600 148836
rect 321000 148336 321100 148736
rect 321500 148336 321600 148736
rect 321000 148236 321600 148336
rect 316358 147826 316414 147836
rect 315854 146701 315910 147470
rect 314090 146576 314146 146616
rect 313838 146454 313894 146494
rect 313586 146332 313642 146372
rect 313334 146210 313390 146250
rect 313082 146088 313138 146128
rect 312830 145966 312886 146006
rect 312578 145844 312634 145884
rect 312326 145722 312382 145762
rect 312074 145600 312130 145640
rect 311822 145478 311878 145518
rect 311570 145356 311626 145396
rect 311318 145234 311374 145274
rect 311066 145112 311122 145152
rect 310814 144990 310870 145030
rect 310562 144868 310618 144908
rect 310310 144746 310366 144786
rect 310058 144624 310114 144664
rect 309806 144502 309862 144542
rect 309554 144380 309610 144420
rect 309302 144258 309358 144298
rect 309050 144136 309106 144176
rect 308798 144014 308854 144054
rect 308546 143892 308602 143932
rect 308294 143770 308350 143810
rect 308042 143648 308098 143688
rect 307790 143526 307846 143566
rect 307538 143404 307594 143444
rect 307286 143282 307342 143322
rect 307034 143160 307090 143200
rect 306782 143038 306838 143078
rect 306530 142916 306586 142956
rect 306278 142794 306334 142834
rect 306026 142672 306082 142712
rect 305774 142550 305830 142590
rect 305522 142428 305578 142468
rect 305270 142306 305326 142346
rect 305018 142184 305074 142224
rect 304766 142062 304822 142102
rect 304514 141940 304570 141980
rect 304262 141818 304318 141858
rect 304010 141696 304066 141736
rect 303758 141574 303814 141614
rect 303506 141452 303562 141492
rect 303254 141330 303310 141370
rect 303002 141208 303058 141248
rect 302750 141086 302806 141126
rect 302498 140964 302554 141004
rect 302246 140842 302302 140882
rect 301994 140720 302050 140760
rect 301742 140598 301798 140638
rect 301490 140476 301546 140516
rect 301238 140354 301294 140394
rect 300986 140232 301042 140272
rect 300734 140110 300790 140150
rect 300482 139988 300538 140028
rect 300230 139866 300286 139906
rect 299978 139744 300034 139784
rect 299726 139622 299782 139662
rect 299474 139500 299530 139540
rect 299222 139378 299278 139418
rect 298970 139256 299026 139296
rect 298718 139134 298774 139174
rect 298466 139012 298522 139052
rect 298214 138890 298270 138930
rect 297962 138768 298018 138808
rect 297710 138646 297766 138686
rect 297458 138524 297514 138564
rect 297206 138402 297262 138442
rect 296954 138280 297010 138320
rect 296702 138158 296758 138198
rect 296450 138036 296506 138076
rect 296198 137914 296254 137954
rect 295694 137766 295750 137798
rect 295946 137792 296002 137832
rect 295694 64654 295750 137710
rect 479150 122610 479206 338232
rect 479150 122448 479206 122488
rect 479402 117242 479458 338476
rect 479654 117852 479710 338720
rect 479906 134566 479962 338964
rect 479906 134404 479962 134444
rect 480158 134078 480214 339208
rect 480410 139446 480466 339452
rect 480662 337516 480718 370514
rect 480662 337420 480718 337460
rect 481908 369376 481964 369488
rect 481670 337272 481726 337326
rect 481418 337028 481474 337082
rect 481166 336784 481222 336838
rect 480914 336540 480970 336594
rect 480914 298046 480970 336484
rect 481166 331596 481222 336728
rect 481166 331434 481222 331474
rect 481418 314882 481474 336972
rect 481418 314720 481474 314760
rect 481670 298656 481726 337216
rect 481670 298494 481726 298534
rect 480914 297884 480970 297924
rect 480410 139284 480466 139324
rect 481908 245392 481964 369264
rect 481908 144816 481964 245280
rect 482160 339676 482216 339692
rect 482160 332192 482216 339620
rect 482160 315392 482216 332080
rect 482160 225008 482216 315280
rect 482160 224850 482216 224896
rect 481908 144256 481964 144704
rect 481908 138208 481964 144144
rect 481376 135058 481472 135076
rect 481376 134566 481472 134952
rect 481376 134416 481472 134444
rect 481690 135062 481812 135116
rect 480158 133916 480214 133956
rect 481380 134078 481476 134114
rect 481380 133626 481476 133956
rect 481380 133504 481476 133520
rect 481690 133638 481812 134934
rect 479654 117690 479710 117730
rect 481376 118258 481472 118276
rect 481376 117852 481472 118152
rect 481376 117702 481472 117730
rect 481690 118262 481812 133510
rect 479402 117080 479458 117120
rect 481380 117242 481476 117278
rect 481380 116826 481476 117120
rect 481380 116704 481476 116720
rect 481690 116838 481812 118134
rect 481690 116472 481812 116710
rect 481908 128016 481964 138096
rect 481908 127456 481964 127904
rect 481908 121408 481964 127344
rect 477200 79400 477800 79500
rect 477200 79000 477300 79400
rect 477700 79000 477800 79400
rect 477200 78900 477800 79000
rect 477200 78400 477800 78500
rect 477200 78000 477300 78400
rect 477700 78000 477800 78400
rect 477200 77900 477800 78000
rect 472400 75600 478000 75800
rect 295694 64598 303750 64654
rect 295442 64346 303498 64402
rect 295190 64094 303246 64150
rect 294938 63842 302994 63898
rect 294686 63590 302742 63646
rect 294434 63338 302490 63394
rect 294182 63086 302238 63142
rect 293930 62834 301986 62890
rect 293678 62582 301734 62638
rect 293426 62330 301482 62386
rect 293174 62078 301230 62134
rect 292922 61826 300978 61882
rect 292670 61574 300726 61630
rect 268380 61362 283248 61488
rect 268380 59472 268506 61362
rect 283122 59472 283248 61362
rect 268380 59346 283248 59472
rect 285200 58600 300000 58800
rect 285200 53400 285400 58600
rect 299800 53400 300000 58600
rect 285200 53200 300000 53400
rect 231600 42200 246400 42400
rect 231600 37200 231800 42200
rect 246200 37200 246400 42200
rect 231600 37000 246400 37200
rect 300670 34980 300726 61574
rect 300922 35164 300978 61826
rect 301174 35408 301230 62078
rect 301426 35652 301482 62330
rect 301678 35896 301734 62582
rect 301930 36140 301986 62834
rect 302182 36384 302238 63086
rect 302434 36628 302490 63338
rect 302686 36872 302742 63590
rect 302938 37116 302994 63842
rect 303190 37360 303246 64094
rect 303442 37604 303498 64346
rect 303694 37848 303750 64598
rect 472400 61200 472600 75600
rect 477800 61200 478000 75600
rect 472400 61000 478000 61200
rect 317800 52300 318600 52400
rect 317800 51700 317900 52300
rect 318500 51700 318600 52300
rect 317800 51600 318600 51700
rect 317800 51100 318600 51200
rect 317800 50500 317900 51100
rect 318500 50500 318600 51100
rect 317800 50400 318600 50500
rect 481418 49044 481474 49072
rect 480400 45100 481200 45200
rect 480400 44500 480500 45100
rect 481100 44500 481200 45100
rect 480400 44400 481200 44500
rect 480400 43700 481200 43800
rect 480400 43100 480500 43700
rect 481100 43100 481200 43700
rect 480400 43000 481200 43100
rect 481418 37848 481474 48922
rect 303694 37792 481474 37848
rect 481908 47824 481964 121296
rect 303442 37548 328104 37604
rect 328230 37548 328270 37604
rect 303190 37304 420714 37360
rect 420840 37304 420880 37360
rect 302938 37060 403956 37116
rect 404082 37060 404122 37116
rect 302686 36816 387072 36872
rect 387198 36816 387238 36872
rect 302434 36572 370314 36628
rect 370440 36572 370480 36628
rect 302182 36328 311346 36384
rect 311472 36328 311512 36384
rect 301930 36084 311976 36140
rect 312102 36084 312142 36140
rect 301678 35840 328734 35896
rect 328860 35840 328900 35896
rect 301426 35596 365526 35652
rect 365652 35596 365692 35652
rect 301174 35352 382284 35408
rect 382410 35352 382450 35408
rect 300922 35108 399168 35164
rect 399294 35108 399334 35164
rect 218234 34913 300244 34969
rect 300300 34913 300310 34969
rect 300670 34924 415926 34980
rect 416052 34924 416092 34980
rect 217520 34630 364896 34686
rect 365022 34630 365148 34686
rect 217268 34378 381654 34434
rect 381780 34378 381906 34434
rect 217016 34126 398538 34182
rect 398664 34126 398790 34182
rect 216764 33874 415296 33930
rect 415422 33874 415462 33930
rect 216512 33606 471492 33662
rect 471618 33606 471744 33662
rect 33054 33372 56538 33428
rect 56594 33372 56634 33428
rect 481908 33404 481964 47712
rect 300234 33348 300244 33404
rect 300300 33348 369040 33404
rect 369152 33348 385840 33404
rect 385952 33348 402640 33404
rect 402752 33348 419440 33404
rect 419552 33348 470288 33404
rect 470400 33348 481964 33404
rect 32802 33120 90180 33176
rect 90236 33120 90276 33176
rect 310648 33078 310886 33200
rect 311014 33078 312310 33200
rect 312438 33078 327686 33200
rect 327814 33078 329110 33200
rect 329238 33078 364486 33200
rect 364614 33078 365910 33200
rect 366038 33078 381286 33200
rect 381414 33078 382710 33200
rect 382838 33078 398086 33200
rect 398214 33078 399510 33200
rect 399638 33078 414886 33200
rect 415014 33078 416310 33200
rect 416438 33078 432820 33200
rect 433812 33078 433869 33200
rect 310880 32768 310896 32864
rect 311002 32768 311346 32864
rect 311472 32768 311504 32864
rect 311952 32764 311976 32860
rect 312102 32764 312328 32860
rect 312434 32764 312452 32860
rect 327680 32768 327696 32864
rect 327802 32768 328104 32864
rect 328230 32768 328262 32864
rect 328710 32764 328734 32860
rect 328860 32764 329128 32860
rect 329234 32764 329252 32860
rect 364480 32768 364496 32864
rect 364602 32768 364896 32864
rect 365022 32768 365054 32864
rect 365502 32764 365526 32860
rect 365652 32764 365928 32860
rect 366034 32764 366052 32860
rect 381280 32768 381296 32864
rect 381402 32768 381654 32864
rect 381780 32768 381812 32864
rect 382260 32764 382284 32860
rect 382410 32764 382728 32860
rect 382834 32764 382852 32860
rect 398080 32768 398096 32864
rect 398202 32768 398538 32864
rect 398664 32768 398696 32864
rect 399144 32764 399168 32860
rect 399294 32764 399528 32860
rect 399634 32764 399652 32860
rect 414880 32768 414896 32864
rect 415002 32768 415296 32864
rect 415422 32768 415454 32864
rect 415902 32764 415926 32860
rect 416052 32764 416328 32860
rect 416434 32764 416452 32860
rect 32550 32624 55404 32680
rect 55460 32624 72162 32680
rect 72218 32624 88920 32680
rect 88976 32624 89016 32680
<< via2 >>
rect 78708 381220 78764 381276
rect 80052 381108 80108 381164
rect 82628 380996 82684 381052
rect 82740 380884 82796 380940
rect 85428 380772 85484 380828
rect 78820 380660 78876 380716
rect 80164 380548 80220 380604
rect 82516 380436 82572 380492
rect 33600 366000 34600 380400
rect 82852 380324 82908 380380
rect 85652 380212 85708 380268
rect 332154 380250 332744 380778
rect 78932 380100 78988 380156
rect 80276 379988 80332 380044
rect 82404 379876 82460 379932
rect 82964 379764 83020 379820
rect 85876 379652 85932 379708
rect 79044 379540 79100 379596
rect 80388 379428 80444 379484
rect 82292 379316 82348 379372
rect 83076 379204 83132 379260
rect 79156 379092 79212 379148
rect 80500 378980 80556 379036
rect 82180 378868 82236 378924
rect 83188 378756 83244 378812
rect 79268 378644 79324 378700
rect 80612 378532 80668 378588
rect 82068 378420 82124 378476
rect 83300 378308 83356 378364
rect 79380 378196 79436 378252
rect 80724 378084 80780 378140
rect 81956 377972 82012 378028
rect 83412 377860 83468 377916
rect 79492 377748 79548 377804
rect 80836 377636 80892 377692
rect 81844 377524 81900 377580
rect 83524 377412 83580 377468
rect 79604 377300 79660 377356
rect 80948 377188 81004 377244
rect 81732 377076 81788 377132
rect 83636 376964 83692 377020
rect 79716 376852 79772 376908
rect 81060 376740 81116 376796
rect 81620 376628 81676 376684
rect 83748 376516 83804 376572
rect 79828 376404 79884 376460
rect 81172 376292 81228 376348
rect 81508 376180 81564 376236
rect 83860 376068 83916 376124
rect 79940 375956 79996 376012
rect 81284 375844 81340 375900
rect 81396 375732 81452 375788
rect 83972 375620 84028 375676
rect 78708 372624 78764 373072
rect 68964 370730 69020 370786
rect 68852 370486 68908 370542
rect 63504 366912 64764 367542
rect 68292 366094 68348 366150
rect 33600 349200 34600 363600
rect 68068 362190 68124 362246
rect 65394 360360 65646 360864
rect 66150 360360 66780 361620
rect 64092 359493 64148 359549
rect 63126 358092 63378 358470
rect 64764 359269 64820 359325
rect 68068 359493 68124 359549
rect 68292 359269 68348 359325
rect 68516 365606 68572 365662
rect 65050 359045 65106 359101
rect 68516 359045 68572 359101
rect 68740 364386 68796 364442
rect 33120 335888 33462 336226
rect 32676 285572 32732 285628
rect 32788 286356 32844 286412
rect 32564 285124 32620 285180
rect 32340 284228 32396 284284
rect 32452 284676 32508 284732
rect 33348 286244 33404 286300
rect 33236 285684 33292 285740
rect 33124 285236 33180 285292
rect 33012 284788 33068 284844
rect 33908 286132 33964 286188
rect 33796 285796 33852 285852
rect 33684 285348 33740 285404
rect 33572 284900 33628 284956
rect 34580 336980 34636 337036
rect 34468 286020 34524 286076
rect 34356 285908 34412 285964
rect 34244 285460 34300 285516
rect 34132 285012 34188 285068
rect 34020 284564 34076 284620
rect 33460 284452 33516 284508
rect 32900 284340 32956 284396
rect 33526 283714 33670 283874
rect 33739 254062 33994 257206
rect 68516 336980 68572 337036
rect 36726 315029 36786 315085
rect 41151 314906 41211 314966
rect 44138 315029 44198 315085
rect 46265 314906 46325 314966
rect 41326 314673 41386 314729
rect 42308 314785 42364 314841
rect 36486 313906 36546 313966
rect 35154 312984 35910 313488
rect 38413 313438 38578 313604
rect 38413 313329 38578 313438
rect 39889 313438 40051 313597
rect 39889 313333 40051 313438
rect 41744 313438 41962 313623
rect 41744 313357 41962 313438
rect 42532 314561 42588 314617
rect 42840 312858 43218 313614
rect 44030 313428 44407 313687
rect 45467 313456 45631 313601
rect 45467 313339 45631 313456
rect 46871 314673 46931 314729
rect 47959 314673 48019 314729
rect 62343 315027 62400 315084
rect 49364 314357 49420 314413
rect 46935 313456 47111 313610
rect 46935 313336 47111 313456
rect 48779 313456 49011 313634
rect 48779 313364 49011 313456
rect 42840 310338 43218 310842
rect 49588 314133 49644 314189
rect 60354 313110 61236 313362
rect 56644 312117 56700 312173
rect 60354 311472 61236 311724
rect 65750 314979 65826 315035
rect 62692 313908 62748 313964
rect 64135 313907 64192 313964
rect 63084 313685 63140 313741
rect 64512 312480 65394 312732
rect 50022 310338 50400 310842
rect 64184 310716 64240 310842
rect 64520 310535 64596 310611
rect 50652 309078 51282 309582
rect 57903 310206 58105 310424
rect 58590 308952 58842 309582
rect 52708 308528 52947 308767
rect 51619 308134 51968 308285
rect 66048 314979 66108 315035
rect 66228 314979 66288 315035
rect 65927 313461 65984 313517
rect 67719 313237 67776 313293
rect 68852 314805 68908 314861
rect 68964 314581 69020 314637
rect 69076 369266 69132 369322
rect 69076 314357 69132 314413
rect 69188 369022 69244 369078
rect 69188 314133 69244 314189
rect 69300 365362 69356 365418
rect 69636 364874 69692 364930
rect 69524 364630 69580 364686
rect 69300 313909 69356 313965
rect 69412 362434 69468 362490
rect 69412 313685 69468 313741
rect 69524 313461 69580 313517
rect 74452 364142 74508 364198
rect 71652 363898 71708 363954
rect 71540 363654 71596 363710
rect 71428 363410 71484 363466
rect 71316 361702 71372 361758
rect 69636 313237 69692 313293
rect 69748 357066 69804 357122
rect 68740 312117 68796 312173
rect 65976 310716 66032 310842
rect 68670 310968 69426 311220
rect 67768 310716 67824 310842
rect 67446 310535 67522 310611
rect 68976 283922 69088 284032
rect 37740 281653 38303 282078
rect 37590 248893 38138 249473
rect 58590 247086 59220 247968
rect 60228 245448 60858 246330
rect 63882 243936 64638 244692
rect 46116 243728 46172 243784
rect 34339 237262 34594 240406
rect 33176 219357 33382 223223
rect 64036 243728 64092 243784
rect 46116 240816 46172 240872
rect 47908 243606 47964 243662
rect 62244 243606 62300 243662
rect 47908 240694 47964 240750
rect 49700 243484 49756 243540
rect 60452 243484 60508 243540
rect 49700 240572 49756 240628
rect 51492 243362 51548 243418
rect 58660 243362 58716 243418
rect 51492 240450 51548 240506
rect 53284 243240 53340 243296
rect 56868 243240 56924 243296
rect 53284 240328 53340 240384
rect 55076 243118 55132 243174
rect 55076 240206 55132 240262
rect 56868 240084 56924 240140
rect 58660 239962 58716 240018
rect 49770 239778 51660 239904
rect 60452 239840 60508 239896
rect 62244 239718 62300 239774
rect 67284 242298 67914 243180
rect 65764 241290 66898 241794
rect 64036 239596 64092 239652
rect 37740 237453 38303 237878
rect 64849 233982 65109 234149
rect 69860 356822 69916 356878
rect 70084 356578 70140 356634
rect 69972 356334 70028 356390
rect 71204 353650 71260 353706
rect 71092 353406 71148 353462
rect 70980 353162 71036 353218
rect 70868 352918 70924 352974
rect 70756 352674 70812 352730
rect 70644 352430 70700 352486
rect 70532 352186 70588 352242
rect 70420 351942 70476 351998
rect 70308 351698 70364 351754
rect 70196 351454 70252 351510
rect 73220 363166 73276 363222
rect 73108 362922 73164 362978
rect 72996 362678 73052 362734
rect 72884 361458 72940 361514
rect 71764 351210 71820 351266
rect 71876 350966 71932 351022
rect 71988 350722 72044 350778
rect 72100 350478 72156 350534
rect 72212 350234 72268 350290
rect 72324 349990 72380 350046
rect 72436 349746 72492 349802
rect 72548 349502 72604 349558
rect 72660 349258 72716 349314
rect 72772 349014 72828 349070
rect 73332 356090 73388 356146
rect 73332 240816 73388 240872
rect 73444 355846 73500 355902
rect 73444 240694 73500 240750
rect 73556 355602 73612 355658
rect 73556 240572 73612 240628
rect 73668 355358 73724 355414
rect 73668 240450 73724 240506
rect 73780 355114 73836 355170
rect 73780 240328 73836 240384
rect 73892 354870 73948 354926
rect 73892 240206 73948 240262
rect 74004 354626 74060 354682
rect 74004 240084 74060 240140
rect 74116 354382 74172 354438
rect 74116 239962 74172 240018
rect 74228 354138 74284 354194
rect 74228 239840 74284 239896
rect 74340 353894 74396 353950
rect 74340 239718 74396 239774
rect 78820 372624 78876 373072
rect 76356 285908 76412 285964
rect 76244 285796 76300 285852
rect 76132 285684 76188 285740
rect 76020 285572 76076 285628
rect 75908 285460 75964 285516
rect 75796 285348 75852 285404
rect 75684 285236 75740 285292
rect 75572 285124 75628 285180
rect 75460 285012 75516 285068
rect 75348 284900 75404 284956
rect 75236 284788 75292 284844
rect 75124 284676 75180 284732
rect 75012 284564 75068 284620
rect 74900 284452 74956 284508
rect 74788 284340 74844 284396
rect 74676 284228 74732 284284
rect 75572 256904 75628 256960
rect 75684 256660 75740 256716
rect 75796 256416 75852 256472
rect 76356 257880 76412 257936
rect 76244 257636 76300 257692
rect 76132 257392 76188 257448
rect 76020 257148 76076 257204
rect 75908 256172 75964 256228
rect 75460 250072 75516 250128
rect 75348 249828 75404 249884
rect 75236 249584 75292 249640
rect 75124 249340 75180 249396
rect 78932 372624 78988 373072
rect 79044 372624 79100 373072
rect 79156 372624 79212 373072
rect 79268 372624 79324 373072
rect 79380 372624 79436 373072
rect 79492 372624 79548 373072
rect 79604 372624 79660 373072
rect 79716 372624 79772 373072
rect 79828 372624 79884 373072
rect 79940 372624 79996 373072
rect 80052 372624 80108 373072
rect 80164 372624 80220 373072
rect 80276 372624 80332 373072
rect 80388 372624 80444 373072
rect 80500 372624 80556 373072
rect 80612 372624 80668 373072
rect 80724 372624 80780 373072
rect 80836 372624 80892 373072
rect 80948 372624 81004 373072
rect 81060 372624 81116 373072
rect 81172 372624 81228 373072
rect 81284 372624 81340 373072
rect 81396 372624 81452 373072
rect 81508 372624 81564 373072
rect 81620 372624 81676 373072
rect 81732 372624 81788 373072
rect 81844 372624 81900 373072
rect 81956 372624 82012 373072
rect 82068 372624 82124 373072
rect 82180 372624 82236 373072
rect 82292 372624 82348 373072
rect 82404 372624 82460 373072
rect 82516 372624 82572 373072
rect 82628 372624 82684 373072
rect 82740 372624 82796 373072
rect 82852 372624 82908 373072
rect 82964 372624 83020 373072
rect 83076 372624 83132 373072
rect 83188 372624 83244 373072
rect 83300 372624 83356 373072
rect 83412 372624 83468 373072
rect 83524 372624 83580 373072
rect 83636 372624 83692 373072
rect 83748 372624 83804 373072
rect 83860 372624 83916 373072
rect 83972 372624 84028 373072
rect 85428 372624 85484 373072
rect 84980 366094 85036 366150
rect 84084 361214 84140 361270
rect 84308 360970 84364 361026
rect 82740 286356 82796 286412
rect 84532 360726 84588 360782
rect 82964 286244 83020 286300
rect 84756 360482 84812 360538
rect 83188 286132 83244 286188
rect 85428 360238 85484 360294
rect 85652 372624 85708 373072
rect 85652 359994 85708 360050
rect 85876 372624 85932 373072
rect 88424 371234 88480 371290
rect 87164 370982 87220 371038
rect 85876 359750 85932 359806
rect 86156 368778 86212 368834
rect 84980 348526 85036 348582
rect 85358 348038 85414 348094
rect 83412 286020 83468 286076
rect 85092 346574 85148 346630
rect 82628 266582 82684 266638
rect 82516 260564 82572 260620
rect 82404 260320 82460 260376
rect 82292 260076 82348 260132
rect 82180 259832 82236 259888
rect 82068 259588 82124 259644
rect 81956 259344 82012 259400
rect 81844 259100 81900 259156
rect 81732 258856 81788 258912
rect 81620 258612 81676 258668
rect 81508 258368 81564 258424
rect 81396 258124 81452 258180
rect 81284 255928 81340 255984
rect 81172 255684 81228 255740
rect 81060 255440 81116 255496
rect 80948 255196 81004 255252
rect 80836 254952 80892 255008
rect 80724 254708 80780 254764
rect 80612 254464 80668 254520
rect 80500 254220 80556 254276
rect 80388 253976 80444 254032
rect 80276 253732 80332 253788
rect 80164 253488 80220 253544
rect 80052 253244 80108 253300
rect 79940 253000 79996 253056
rect 79828 252756 79884 252812
rect 79716 252512 79772 252568
rect 79604 252268 79660 252324
rect 79492 252024 79548 252080
rect 79380 251780 79436 251836
rect 79268 251536 79324 251592
rect 79156 251292 79212 251348
rect 79044 251048 79100 251104
rect 78932 250804 78988 250860
rect 78820 250560 78876 250616
rect 78708 250316 78764 250372
rect 78596 249096 78652 249152
rect 78484 248852 78540 248908
rect 78372 248608 78428 248664
rect 78260 248364 78316 248420
rect 78148 248120 78204 248176
rect 78036 247876 78092 247932
rect 77924 247632 77980 247688
rect 77812 247388 77868 247444
rect 77700 247144 77756 247200
rect 77588 246900 77644 246956
rect 77476 246656 77532 246712
rect 77364 246412 77420 246468
rect 75012 246168 75068 246224
rect 74900 245924 74956 245980
rect 74788 245680 74844 245736
rect 74676 245436 74732 245492
rect 74452 239596 74508 239652
rect 66402 232596 66654 233604
rect 64234 225689 64745 226767
rect 72450 228690 73584 229320
rect 72954 208656 73584 209538
rect 34939 203662 35194 206806
rect 35539 186862 35794 190006
rect 79331 206980 79685 207942
rect 73444 206658 73500 206714
rect 37590 205293 38138 205873
rect 74116 206546 74172 206602
rect 73780 205944 73836 206000
rect 73780 203268 73836 203324
rect 74788 206434 74844 206490
rect 74345 205038 74614 205722
rect 75460 206322 75516 206378
rect 75124 205944 75180 206000
rect 75124 205202 75180 205258
rect 76132 206210 76188 206266
rect 75572 205314 75628 205370
rect 75572 203390 75628 203446
rect 76804 206098 76860 206154
rect 77476 205986 77532 206042
rect 77364 205426 77420 205482
rect 77364 203512 77420 203568
rect 78148 205874 78204 205930
rect 78820 205762 78876 205818
rect 79492 205650 79548 205706
rect 79492 203146 79548 203202
rect 78820 203024 78876 203080
rect 78148 202902 78204 202958
rect 77476 202780 77532 202836
rect 76804 202658 76860 202714
rect 76132 202536 76188 202592
rect 75460 202414 75516 202470
rect 74788 202292 74844 202348
rect 74116 202170 74172 202226
rect 73444 202048 73500 202104
rect 73206 199710 73710 200970
rect 64545 198151 64831 198350
rect 49829 196869 51830 197117
rect 37740 194653 38303 195078
rect 70812 198094 71316 198850
rect 65443 197377 65722 197670
rect 69048 192402 69552 193032
rect 80164 205538 80220 205594
rect 80164 203634 80220 203690
rect 66150 189252 66780 190008
rect 64260 182952 64764 184338
rect 66801 185801 67014 185968
rect 67014 185801 67096 185968
rect 36139 170062 36394 173206
rect 36739 153262 36994 156406
rect 32998 146020 33054 146076
rect 32550 122368 32606 122424
rect 32550 118958 32606 119202
rect 32802 145760 32858 145816
rect 73332 166446 74088 167202
rect 79506 164178 79884 165312
rect 73444 163836 73500 163892
rect 37590 162493 38138 163073
rect 80388 163836 80444 163892
rect 74116 163724 74172 163780
rect 73780 162380 73836 162436
rect 73780 160446 73836 160502
rect 80500 163724 80556 163780
rect 74788 163612 74844 163668
rect 80612 163612 80668 163668
rect 75460 163500 75516 163556
rect 80724 163500 80780 163556
rect 76132 163388 76188 163444
rect 75572 162492 75628 162548
rect 75572 160568 75628 160624
rect 80836 163388 80892 163444
rect 76804 163276 76860 163332
rect 80948 163276 81004 163332
rect 77476 163164 77532 163220
rect 77364 162604 77420 162660
rect 77364 160690 77420 160746
rect 81060 163164 81116 163220
rect 78148 163052 78204 163108
rect 81172 163052 81228 163108
rect 78820 162940 78876 162996
rect 81284 162940 81340 162996
rect 79492 162828 79548 162884
rect 81396 162828 81452 162884
rect 80164 162716 80220 162772
rect 81508 162716 81564 162772
rect 81620 162604 81676 162660
rect 81732 162492 81788 162548
rect 81956 206658 82012 206714
rect 82068 206546 82124 206602
rect 82180 206434 82236 206490
rect 82292 206322 82348 206378
rect 82404 206210 82460 206266
rect 82516 206098 82572 206154
rect 82628 205986 82684 206042
rect 82740 205874 82796 205930
rect 82852 205762 82908 205818
rect 82964 205650 83020 205706
rect 83076 205538 83132 205594
rect 83188 205426 83244 205482
rect 83300 205314 83356 205370
rect 83412 205202 83468 205258
rect 81844 162380 81900 162436
rect 80892 161532 81522 162036
rect 80164 160812 80220 160868
rect 79492 160324 79548 160380
rect 78820 160202 78876 160258
rect 78148 160080 78204 160136
rect 77476 159958 77532 160014
rect 76804 159836 76860 159892
rect 76132 159714 76188 159770
rect 75460 159592 75516 159648
rect 74788 159470 74844 159526
rect 74116 159348 74172 159404
rect 73444 159226 73500 159282
rect 70964 156500 71720 156752
rect 72072 156492 72828 156744
rect 61684 155540 61740 155596
rect 60004 155400 60060 155456
rect 51408 152838 52794 153468
rect 37156 146020 37212 146076
rect 47236 145908 47292 145964
rect 52500 146580 52556 146636
rect 53060 146356 53116 146412
rect 53620 146132 53676 146188
rect 54180 145908 54236 145964
rect 55524 146132 55580 146188
rect 56644 146356 56700 146412
rect 56868 146580 56924 146636
rect 32998 143556 33054 143612
rect 32802 143332 32858 143388
rect 32802 118958 32858 119202
rect 33054 143108 33110 143164
rect 33054 118958 33110 119202
rect 33306 142884 33362 142940
rect 33306 118958 33362 119202
rect 33558 142660 33614 142716
rect 33558 118958 33614 119202
rect 33810 142436 33866 142492
rect 58548 139972 58604 140028
rect 58324 137284 58380 137340
rect 52276 123508 52332 123564
rect 52500 123732 52556 123788
rect 52724 123956 52780 124012
rect 53284 124180 53340 124236
rect 56308 124404 56364 124460
rect 52052 123284 52108 123340
rect 51828 123060 51884 123116
rect 48916 122836 48972 122892
rect 44324 122612 44380 122668
rect 39360 121492 39428 121548
rect 39232 121268 39300 121324
rect 39104 121044 39172 121100
rect 33810 118958 33866 119202
rect 38976 120820 39044 120876
rect 34650 114912 35406 116046
rect 34333 101246 34506 109085
rect 37674 108612 38556 109620
rect 37870 107984 38167 108040
rect 37870 107648 38167 107704
rect 61796 155278 61852 155334
rect 61334 143810 61390 143866
rect 62356 155156 62412 155212
rect 62468 155034 62524 155090
rect 61908 139076 61964 139132
rect 63028 154912 63084 154968
rect 63140 154790 63196 154846
rect 62580 138852 62636 138908
rect 63700 154668 63756 154724
rect 63812 154546 63868 154602
rect 63252 138628 63308 138684
rect 64372 154424 64428 154480
rect 64484 154302 64540 154358
rect 63924 138404 63980 138460
rect 60984 133560 61362 135828
rect 65044 154180 65100 154236
rect 65156 154058 65212 154114
rect 64596 138180 64652 138236
rect 65716 153936 65772 153992
rect 65828 153814 65884 153870
rect 65268 137956 65324 138012
rect 66388 153692 66444 153748
rect 66500 153570 66556 153626
rect 65940 137732 65996 137788
rect 67060 153448 67116 153504
rect 67172 153326 67228 153382
rect 66612 137508 66668 137564
rect 67732 153204 67788 153260
rect 67844 153082 67900 153138
rect 67284 142660 67340 142716
rect 68404 152838 68460 152894
rect 68850 152716 68910 152772
rect 67956 142436 68012 142492
rect 68628 142212 68684 142268
rect 69076 152594 69132 152650
rect 69636 152472 69692 152528
rect 69300 141988 69356 142044
rect 66612 131908 66668 131964
rect 62748 131040 65646 131292
rect 59875 130503 60078 130511
rect 59875 130447 60078 130503
rect 59875 130057 60078 130447
rect 61634 130445 61874 130477
rect 61634 130051 61874 130445
rect 62748 130158 65646 130410
rect 60340 127988 60396 128044
rect 59850 127386 60102 127638
rect 61110 126630 61866 127008
rect 59114 124628 59194 124684
rect 67172 131908 67228 131964
rect 69748 152350 69804 152406
rect 70308 152228 70364 152284
rect 69972 141764 70028 141820
rect 67732 131908 67788 131964
rect 68852 131908 68908 131964
rect 68964 130577 69020 130633
rect 68964 128884 69020 128940
rect 70420 152106 70476 152162
rect 70980 151984 71036 152040
rect 70644 141540 70700 141596
rect 69412 131908 69468 131964
rect 70532 136276 70588 136332
rect 71092 151862 71148 151918
rect 71652 151740 71708 151796
rect 71316 141316 71372 141372
rect 71204 136052 71260 136108
rect 71764 151618 71820 151674
rect 72324 151496 72380 151552
rect 71988 141092 72044 141148
rect 69972 131908 70028 131964
rect 70532 131908 70588 131964
rect 69860 129780 69916 129836
rect 69188 128212 69244 128268
rect 67396 126196 67452 126252
rect 66612 124852 66668 124908
rect 66612 122368 66668 122424
rect 70550 121716 70606 121772
rect 58324 107984 58380 108040
rect 59000 110054 59056 110110
rect 39560 106453 39628 106605
rect 41220 106254 41288 106310
rect 70980 110054 71036 110110
rect 72436 151374 72492 151430
rect 72996 151252 73052 151308
rect 72660 140868 72716 140924
rect 66906 108738 67536 109116
rect 61486 107648 61546 107704
rect 59598 106974 60606 107352
rect 71008 108500 71450 108556
rect 65898 107226 66528 107604
rect 59000 106254 59056 106310
rect 62384 106198 62658 106254
rect 72548 137284 72604 137340
rect 73108 151130 73164 151186
rect 73668 151008 73724 151064
rect 73332 140644 73388 140700
rect 73220 137060 73276 137116
rect 73780 150886 73836 150942
rect 74340 150764 74396 150820
rect 74004 140420 74060 140476
rect 74452 150642 74508 150698
rect 75012 150520 75068 150576
rect 74676 140196 74732 140252
rect 72314 132174 73070 132804
rect 71876 131572 71932 131628
rect 73892 124404 73948 124460
rect 75124 150398 75180 150454
rect 75684 150276 75740 150332
rect 75348 143556 75404 143612
rect 74564 124180 74620 124236
rect 75796 150154 75852 150210
rect 76356 150032 76412 150088
rect 76020 143332 76076 143388
rect 74340 121492 74396 121548
rect 75236 123956 75292 124012
rect 76468 149910 76524 149966
rect 77028 149788 77084 149844
rect 76692 143108 76748 143164
rect 75012 121268 75068 121324
rect 75908 123732 75964 123788
rect 77140 149666 77196 149722
rect 77812 149544 77868 149600
rect 78484 149422 78540 149478
rect 79156 149300 79212 149356
rect 79828 149178 79884 149234
rect 77364 142884 77420 142940
rect 78036 139748 78092 139804
rect 78708 139524 78764 139580
rect 80500 148080 80556 148136
rect 79380 139300 79436 139356
rect 75684 121044 75740 121100
rect 77252 123508 77308 123564
rect 76580 122612 76636 122668
rect 77924 123284 77980 123340
rect 78596 123060 78652 123116
rect 79268 122836 79324 122892
rect 79716 122612 79772 122668
rect 79044 122388 79100 122444
rect 78372 122164 78428 122220
rect 77700 121940 77756 121996
rect 80500 121716 80556 121772
rect 80836 147836 80892 147892
rect 76356 120820 76412 120876
rect 81270 142380 81648 146412
rect 82494 144633 83152 144978
rect 83748 155540 83804 155596
rect 83888 197286 83944 197342
rect 83888 155400 83944 155456
rect 86030 316562 86086 316618
rect 85778 316318 85834 316374
rect 85526 316074 85582 316130
rect 85274 315830 85330 315886
rect 85022 315586 85078 315642
rect 84770 315342 84826 315398
rect 84518 315098 84574 315154
rect 84266 314854 84322 314910
rect 84014 155278 84070 155334
rect 84140 305582 84196 305638
rect 84140 155156 84196 155212
rect 84266 155034 84322 155090
rect 84392 313146 84448 313202
rect 84392 154912 84448 154968
rect 84518 154790 84574 154846
rect 84644 313390 84700 313446
rect 84644 154668 84700 154724
rect 84770 154546 84826 154602
rect 84896 313634 84952 313690
rect 84896 154424 84952 154480
rect 85022 154302 85078 154358
rect 85148 313878 85204 313934
rect 85148 154180 85204 154236
rect 85274 154058 85330 154114
rect 85400 314122 85456 314178
rect 85400 153936 85456 153992
rect 85526 153814 85582 153870
rect 85652 314366 85708 314422
rect 85652 153692 85708 153748
rect 85778 153570 85834 153626
rect 85904 314610 85960 314666
rect 85904 153448 85960 153504
rect 86030 153326 86086 153382
rect 86534 368534 86590 368590
rect 86408 348282 86464 348338
rect 86156 153204 86212 153260
rect 86282 317782 86338 317838
rect 86282 153082 86338 153138
rect 86156 152960 86212 153016
rect 84870 147588 84926 147644
rect 84422 146916 84478 146972
rect 86786 368290 86842 368346
rect 86534 152838 86590 152894
rect 86660 347550 86716 347606
rect 86660 152716 86716 152772
rect 87038 368046 87094 368102
rect 86786 152594 86842 152650
rect 86912 348770 86968 348826
rect 86912 152472 86968 152528
rect 87164 152960 87220 153016
rect 87290 367802 87346 367858
rect 87038 152350 87094 152406
rect 87164 152228 87220 152284
rect 86156 147588 86212 147644
rect 85990 147364 86046 147420
rect 85318 146916 85374 146972
rect 86662 147140 86718 147196
rect 83636 137312 83692 137368
rect 87542 367558 87598 367614
rect 87290 152106 87346 152162
rect 87416 347062 87472 347118
rect 87416 151984 87472 152040
rect 87794 367314 87850 367370
rect 87542 151862 87598 151918
rect 87668 347306 87724 347362
rect 87668 151740 87724 151796
rect 88046 367070 88102 367126
rect 87794 151618 87850 151674
rect 87920 346818 87976 346874
rect 87920 151496 87976 151552
rect 88298 366826 88354 366882
rect 88046 151374 88102 151430
rect 88172 347794 88228 347850
rect 88172 151252 88228 151308
rect 88298 151130 88354 151186
rect 88046 151008 88102 151064
rect 87164 147592 87220 147648
rect 88676 370242 88732 370298
rect 88550 366582 88606 366638
rect 88550 150886 88606 150942
rect 88928 369998 88984 370054
rect 88676 150764 88732 150820
rect 88802 366338 88858 366394
rect 88802 150642 88858 150698
rect 89180 369754 89236 369810
rect 88928 150520 88984 150576
rect 89054 366094 89110 366150
rect 89054 150398 89110 150454
rect 89432 369510 89488 369566
rect 89180 150276 89236 150332
rect 89306 317538 89362 317594
rect 89306 150154 89362 150210
rect 90468 365118 90524 365174
rect 89824 356090 90170 356146
rect 89824 355846 90170 355902
rect 89824 355602 90170 355658
rect 89824 355358 90170 355414
rect 89824 355114 90170 355170
rect 89824 354870 90170 354926
rect 89824 354626 90170 354682
rect 89824 354382 90170 354438
rect 89824 354138 90170 354194
rect 89824 353894 90170 353950
rect 89432 150032 89488 150088
rect 89558 317294 89614 317350
rect 89558 149910 89614 149966
rect 89810 317050 89866 317106
rect 89684 149788 89740 149844
rect 89810 149666 89866 149722
rect 89936 316806 89992 316862
rect 90188 198628 90244 198684
rect 89936 149544 89992 149600
rect 90062 198384 90118 198440
rect 90062 149422 90118 149478
rect 90188 149300 90244 149356
rect 90314 198140 90370 198196
rect 90314 149178 90370 149234
rect 89684 147714 89740 147770
rect 93380 359506 93436 359562
rect 110180 359262 110236 359318
rect 126980 359018 127036 359074
rect 143780 358774 143836 358830
rect 199304 370730 199360 370786
rect 200580 358530 200636 358586
rect 206864 370486 206920 370542
rect 209258 370242 209314 370298
rect 217380 358286 217436 358342
rect 229796 369998 229852 370054
rect 230048 369754 230104 369810
rect 232694 369510 232750 369566
rect 232946 369266 233002 369322
rect 233198 369022 233254 369078
rect 241514 368778 241570 368834
rect 244180 358042 244236 358098
rect 260980 357798 261036 357854
rect 266966 368534 267022 368590
rect 268352 368290 268408 368346
rect 268100 365850 268156 365906
rect 268100 361945 268156 362001
rect 268604 368046 268660 368102
rect 268856 367802 268912 367858
rect 269108 367558 269164 367614
rect 269360 367314 269416 367370
rect 269612 367070 269668 367126
rect 269864 366826 269920 366882
rect 270116 366582 270172 366638
rect 270368 366338 270424 366394
rect 270620 366094 270676 366150
rect 270872 365850 270928 365906
rect 271124 365606 271180 365662
rect 271376 365362 271432 365418
rect 271628 365118 271684 365174
rect 271880 364874 271936 364930
rect 272132 364630 272188 364686
rect 272384 364386 272440 364442
rect 272636 364142 272692 364198
rect 272888 363898 272944 363954
rect 273140 363654 273196 363710
rect 273392 363410 273448 363466
rect 273644 363166 273700 363222
rect 273896 362922 273952 362978
rect 274148 362678 274204 362734
rect 274400 362434 274456 362490
rect 274904 362434 274960 362490
rect 274652 362190 274708 362246
rect 275156 361702 275212 361758
rect 275408 361458 275464 361514
rect 427400 374200 441800 375800
rect 444200 374200 458600 375800
rect 467000 374200 481400 375800
rect 470300 373345 470800 373500
rect 470300 373083 470383 373345
rect 470383 373083 470645 373345
rect 470645 373083 470800 373345
rect 470300 373000 470800 373083
rect 471500 373000 472000 373500
rect 320796 364604 322686 365486
rect 328600 365245 329200 365400
rect 328600 364983 328783 365245
rect 328783 364983 329045 365245
rect 329045 364983 329200 365245
rect 328600 364800 329200 364983
rect 319645 363544 319701 363600
rect 277780 357554 277836 357610
rect 292040 362678 292096 362734
rect 292292 362434 292348 362490
rect 309302 362190 309358 362246
rect 309554 361946 309610 362002
rect 309806 361702 309862 361758
rect 310058 361458 310114 361514
rect 320684 363320 320740 363376
rect 328600 363400 329200 364000
rect 310310 361214 310366 361270
rect 310562 360970 310618 361026
rect 310814 360726 310870 360782
rect 316890 360612 317646 360990
rect 311066 360482 311122 360538
rect 311318 360238 311374 360294
rect 311570 359994 311626 360050
rect 311822 359750 311878 359806
rect 312074 359506 312130 359562
rect 312326 359262 312382 359318
rect 312578 359018 312634 359074
rect 312830 358774 312886 358830
rect 313082 358530 313138 358586
rect 313334 358286 313390 358342
rect 313586 358042 313642 358098
rect 313838 357798 313894 357854
rect 314090 357554 314146 357610
rect 314342 359018 314398 359074
rect 314594 358774 314650 358830
rect 314846 358530 314902 358586
rect 315098 358286 315154 358342
rect 315350 358042 315406 358098
rect 315602 357798 315658 357854
rect 322056 361872 323316 362502
rect 334600 360800 346000 362200
rect 315854 357554 315910 357610
rect 472600 349200 477800 363600
rect 410640 342380 410700 342436
rect 410800 342254 410860 342310
rect 410256 340578 411894 341712
rect 396116 339620 396172 339676
rect 389438 332300 389494 332356
rect 385658 332056 385714 332112
rect 381878 331812 381934 331868
rect 378098 331568 378154 331624
rect 374318 331324 374374 331380
rect 370538 331080 370594 331136
rect 366758 330836 366814 330892
rect 363104 330592 363160 330648
rect 359324 330348 359380 330404
rect 355544 330104 355600 330160
rect 351764 329860 351820 329916
rect 347984 329616 348040 329672
rect 344204 329372 344260 329428
rect 340424 329128 340480 329184
rect 336644 328884 336700 328940
rect 332990 328640 333046 328696
rect 316358 316615 316414 316798
rect 333368 327664 333424 327720
rect 333872 324492 333928 324548
rect 337148 327664 337204 327720
rect 337652 324248 337708 324304
rect 340928 327664 340984 327720
rect 341432 324004 341488 324060
rect 344708 327664 344764 327720
rect 345212 323760 345268 323816
rect 348488 327664 348544 327720
rect 348992 323516 349048 323572
rect 352268 327664 352324 327720
rect 352772 323272 352828 323328
rect 356048 327664 356104 327720
rect 356552 323028 356608 323084
rect 359828 327664 359884 327720
rect 360332 322784 360388 322840
rect 363608 327908 363664 327964
rect 364112 322540 364168 322596
rect 367262 327908 367318 327964
rect 367766 322296 367822 322352
rect 371042 327908 371098 327964
rect 371546 322052 371602 322108
rect 374822 327908 374878 327964
rect 375326 321808 375382 321864
rect 378602 327908 378658 327964
rect 379106 321564 379162 321620
rect 382382 327908 382438 327964
rect 382886 321320 382942 321376
rect 386162 327908 386218 327964
rect 386666 321076 386722 321132
rect 389942 327908 389998 327964
rect 390446 320832 390502 320888
rect 465290 336204 465346 336260
rect 461510 335960 461566 336016
rect 457730 335716 457786 335772
rect 454076 335472 454132 335528
rect 450296 335228 450352 335284
rect 446516 334984 446572 335040
rect 442736 334740 442792 334796
rect 438956 334496 439012 334552
rect 435176 334252 435232 334308
rect 431396 334008 431452 334064
rect 427616 333764 427672 333820
rect 423962 333520 424018 333576
rect 420182 333276 420238 333332
rect 416402 333032 416458 333088
rect 412622 332788 412678 332844
rect 408842 332544 408898 332600
rect 404558 327420 404614 327476
rect 404054 327176 404110 327232
rect 401534 326932 401590 326988
rect 395558 316684 395612 316740
rect 395612 316684 395668 316740
rect 395668 316684 395714 316740
rect 396872 326688 396928 326744
rect 398006 326444 398062 326500
rect 402542 326200 402598 326256
rect 402038 325956 402094 326012
rect 403046 325712 403102 325768
rect 403550 325468 403606 325524
rect 405062 325224 405118 325280
rect 405566 324980 405622 325036
rect 406070 324736 406126 324792
rect 409346 328152 409402 328208
rect 409850 320588 409906 320644
rect 413126 328152 413182 328208
rect 413630 320344 413686 320400
rect 416906 328152 416962 328208
rect 417410 320100 417466 320156
rect 420686 328152 420742 328208
rect 421190 319856 421246 319912
rect 424466 328152 424522 328208
rect 424970 319612 425026 319668
rect 428120 328152 428176 328208
rect 428624 319368 428680 319424
rect 431900 328152 431956 328208
rect 432404 319124 432460 319180
rect 435680 328152 435736 328208
rect 436184 318880 436240 318936
rect 439460 328396 439516 328452
rect 439964 318636 440020 318692
rect 443240 328396 443296 328452
rect 443744 318392 443800 318448
rect 447020 328396 447076 328452
rect 447524 318148 447580 318204
rect 450800 328396 450856 328452
rect 451304 317904 451360 317960
rect 454580 328396 454636 328452
rect 455084 317660 455140 317716
rect 458234 328396 458290 328452
rect 458738 317416 458794 317472
rect 462014 328396 462070 328452
rect 462518 317172 462574 317228
rect 480410 339452 480466 339508
rect 480158 339208 480214 339264
rect 479906 338964 479962 339020
rect 479654 338720 479710 338776
rect 479402 338476 479458 338532
rect 479150 338232 479206 338288
rect 478898 337948 478954 338004
rect 465794 328396 465850 328452
rect 466298 316928 466354 316984
rect 201194 147592 201250 147648
rect 90468 147476 90524 147532
rect 115668 147476 115724 147532
rect 88424 147364 88480 147420
rect 86968 137710 87024 137766
rect 86282 130577 86338 130633
rect 89264 138432 90720 139328
rect 126644 147470 126700 147526
rect 117012 147252 117068 147308
rect 116787 147028 116843 147084
rect 115220 123396 115276 123452
rect 90468 110502 90846 110880
rect 115387 123161 115443 123217
rect 115892 138198 115948 138254
rect 116116 138076 116172 138132
rect 116564 137954 116620 138010
rect 116340 137832 116396 137888
rect 80836 108500 80892 108556
rect 86412 109368 86640 109620
rect 74340 107352 75096 107856
rect 91476 108738 91728 109620
rect 92484 107352 92988 107856
rect 73472 106690 73528 106746
rect 77864 106755 77932 106907
rect 68450 106198 68678 106254
rect 71652 106248 71708 106304
rect 77696 106248 77764 106304
rect 102081 106755 102141 106907
rect 102481 106755 102541 106907
rect 102281 106453 102341 106605
rect 102681 106453 102741 106605
rect 103100 106452 103156 106508
rect 115668 77956 115724 78012
rect 32550 75374 32606 75674
rect 32802 75374 32858 75674
rect 33054 75374 33110 75674
rect 33306 75374 33362 75674
rect 33558 75374 33614 75674
rect 33810 75374 33866 75674
rect 115668 75348 115724 75404
rect 115849 74693 115905 74749
rect 112494 71588 112570 71868
rect 113274 71442 113904 72072
rect 114660 71694 115164 72198
rect 116340 81876 116396 81932
rect 116564 80644 116620 80700
rect 117460 143566 117516 143622
rect 117236 138320 117292 138376
rect 117684 143444 117740 143500
rect 117908 143322 117964 143378
rect 118132 143200 118188 143256
rect 118356 143078 118412 143134
rect 118132 118612 118188 118668
rect 117908 118388 117964 118444
rect 117684 118164 117740 118220
rect 117460 117940 117516 117996
rect 118580 142956 118636 143012
rect 118804 142834 118860 142890
rect 119028 142712 119084 142768
rect 125524 138686 125580 138742
rect 123620 138564 123676 138620
rect 124628 137312 124684 137368
rect 125860 138442 125916 138498
rect 128884 147348 128940 147404
rect 126980 142590 127036 142646
rect 131124 147226 131180 147282
rect 129220 142468 129276 142524
rect 133364 147104 133420 147160
rect 131460 142346 131516 142402
rect 135604 146982 135660 147038
rect 133700 142224 133756 142280
rect 137844 146860 137900 146916
rect 135940 142102 135996 142158
rect 140084 146738 140140 146794
rect 138180 141980 138236 142036
rect 142324 146616 142380 146672
rect 140420 141858 140476 141914
rect 145012 146494 145068 146550
rect 142660 141736 142716 141792
rect 147252 146372 147308 146428
rect 145348 141614 145404 141670
rect 149492 146250 149548 146306
rect 147588 141492 147644 141548
rect 151732 146128 151788 146184
rect 149828 141370 149884 141426
rect 153972 146006 154028 146062
rect 152068 141248 152124 141304
rect 156212 145884 156268 145940
rect 154308 141126 154364 141182
rect 158452 145762 158508 145818
rect 156548 141004 156604 141060
rect 160692 145640 160748 145696
rect 158788 140882 158844 140938
rect 163380 145518 163436 145574
rect 161028 140760 161084 140816
rect 165620 145396 165676 145452
rect 163716 140638 163772 140694
rect 167860 145274 167916 145330
rect 165956 140516 166012 140572
rect 170100 145152 170156 145208
rect 168196 140394 168252 140450
rect 172340 145030 172396 145086
rect 170436 140272 170492 140328
rect 174580 144908 174636 144964
rect 172676 140150 172732 140206
rect 176820 144786 176876 144842
rect 174916 140028 174972 140084
rect 179060 144664 179116 144720
rect 177156 139906 177212 139962
rect 181748 144542 181804 144598
rect 179396 139784 179452 139840
rect 183988 144420 184044 144476
rect 182084 139662 182140 139718
rect 186228 144298 186284 144354
rect 184324 139540 184380 139596
rect 188468 144176 188524 144232
rect 186564 139418 186620 139474
rect 190708 144054 190764 144110
rect 188804 139296 188860 139352
rect 192948 143932 193004 143988
rect 191044 139174 191100 139230
rect 195188 143810 195244 143866
rect 193284 139052 193340 139108
rect 197428 143688 197484 143744
rect 195524 138930 195580 138986
rect 197764 138808 197820 138864
rect 202580 147836 202636 147892
rect 202832 148080 202888 148136
rect 202328 129086 202384 129379
rect 203084 129075 203140 129380
rect 203336 129062 203392 129385
rect 203588 129064 203644 129372
rect 214172 148202 214228 148258
rect 233610 147958 233666 148014
rect 292670 148202 292726 148258
rect 203840 129061 203896 129370
rect 206990 137312 207046 137368
rect 275900 133100 276500 133700
rect 275900 132087 276500 132300
rect 275900 131825 276069 132087
rect 276069 131825 276331 132087
rect 276331 131825 276500 132087
rect 275900 131700 276500 131825
rect 206990 119700 207046 120204
rect 202328 78126 202384 78411
rect 122388 75348 122444 75404
rect 124404 75348 124460 75404
rect 128436 75348 128492 75404
rect 126420 74693 126476 74749
rect 136072 71442 140860 72828
rect 34600 43200 36200 57600
rect 203084 78128 203140 78404
rect 203336 78128 203392 78404
rect 203588 78128 203644 78404
rect 203840 78128 203896 78404
rect 206990 78120 207046 78624
rect 207589 75348 207645 75404
rect 208656 61712 208801 61768
rect 213764 58998 213886 59885
rect 199200 51600 204464 53800
rect 205440 51600 210800 53800
rect 59800 41100 60400 41700
rect 59800 40345 60400 40500
rect 59800 40083 59983 40345
rect 59983 40083 60245 40345
rect 60245 40083 60400 40345
rect 59800 39900 60400 40083
rect 102400 33800 116800 35400
rect 292922 147958 292978 148014
rect 295694 147714 295750 147770
rect 314342 146738 314398 146794
rect 314594 146860 314650 146916
rect 314846 146982 314902 147038
rect 315098 147104 315154 147160
rect 315350 147226 315406 147282
rect 315602 147348 315658 147404
rect 478646 337704 478702 337760
rect 321100 149336 321500 149736
rect 321100 148653 321500 148736
rect 321100 148391 321183 148653
rect 321183 148391 321445 148653
rect 321445 148391 321500 148653
rect 321100 148336 321500 148391
rect 316358 147836 316414 147892
rect 315854 147470 315910 147526
rect 314090 146616 314146 146672
rect 313838 146494 313894 146550
rect 313586 146372 313642 146428
rect 313334 146250 313390 146306
rect 313082 146128 313138 146184
rect 312830 146006 312886 146062
rect 312578 145884 312634 145940
rect 312326 145762 312382 145818
rect 312074 145640 312130 145696
rect 311822 145518 311878 145574
rect 311570 145396 311626 145452
rect 311318 145274 311374 145330
rect 311066 145152 311122 145208
rect 310814 145030 310870 145086
rect 310562 144908 310618 144964
rect 310310 144786 310366 144842
rect 310058 144664 310114 144720
rect 309806 144542 309862 144598
rect 309554 144420 309610 144476
rect 309302 144298 309358 144354
rect 309050 144176 309106 144232
rect 308798 144054 308854 144110
rect 308546 143932 308602 143988
rect 308294 143810 308350 143866
rect 308042 143688 308098 143744
rect 307790 143566 307846 143622
rect 307538 143444 307594 143500
rect 307286 143322 307342 143378
rect 307034 143200 307090 143256
rect 306782 143078 306838 143134
rect 306530 142956 306586 143012
rect 306278 142834 306334 142890
rect 306026 142712 306082 142768
rect 305774 142590 305830 142646
rect 305522 142468 305578 142524
rect 305270 142346 305326 142402
rect 305018 142224 305074 142280
rect 304766 142102 304822 142158
rect 304514 141980 304570 142036
rect 304262 141858 304318 141914
rect 304010 141736 304066 141792
rect 303758 141614 303814 141670
rect 303506 141492 303562 141548
rect 303254 141370 303310 141426
rect 303002 141248 303058 141304
rect 302750 141126 302806 141182
rect 302498 141004 302554 141060
rect 302246 140882 302302 140938
rect 301994 140760 302050 140816
rect 301742 140638 301798 140694
rect 301490 140516 301546 140572
rect 301238 140394 301294 140450
rect 300986 140272 301042 140328
rect 300734 140150 300790 140206
rect 300482 140028 300538 140084
rect 300230 139906 300286 139962
rect 299978 139784 300034 139840
rect 299726 139662 299782 139718
rect 299474 139540 299530 139596
rect 299222 139418 299278 139474
rect 298970 139296 299026 139352
rect 298718 139174 298774 139230
rect 298466 139052 298522 139108
rect 298214 138930 298270 138986
rect 297962 138808 298018 138864
rect 297710 138686 297766 138742
rect 297458 138564 297514 138620
rect 297206 138442 297262 138498
rect 296954 138320 297010 138376
rect 296702 138198 296758 138254
rect 296450 138076 296506 138132
rect 296198 137954 296254 138010
rect 295946 137832 296002 137888
rect 295694 137710 295750 137766
rect 480662 337460 480718 337516
rect 481670 337216 481726 337272
rect 481418 336972 481474 337028
rect 481166 336728 481222 336784
rect 480914 336484 480970 336540
rect 482160 339620 482216 339676
rect 477300 79345 477700 79400
rect 477300 79083 477383 79345
rect 477383 79083 477645 79345
rect 477645 79083 477700 79345
rect 477300 79000 477700 79083
rect 477300 78000 477700 78400
rect 268506 59472 283122 61362
rect 285400 53400 299800 58600
rect 231800 37200 246200 42200
rect 472600 61200 477800 75600
rect 317900 52145 318500 52300
rect 317900 51883 318083 52145
rect 318083 51883 318345 52145
rect 318345 51883 318500 52145
rect 317900 51700 318500 51883
rect 317900 50500 318500 51100
rect 480500 44945 481100 45100
rect 480500 44683 480683 44945
rect 480683 44683 480945 44945
rect 480945 44683 481100 44945
rect 480500 44500 481100 44683
rect 480500 43100 481100 43700
rect 300244 34913 300300 34969
rect 300244 33348 300300 33404
<< metal3 >>
rect 78708 381276 78764 381316
rect 33400 380400 34800 380600
rect 33400 366000 33600 380400
rect 34600 366000 34800 380400
rect 78708 373072 78764 381220
rect 80052 381164 80108 381204
rect 78708 372596 78764 372624
rect 78820 380716 78876 380756
rect 78820 373072 78876 380660
rect 78820 372596 78876 372624
rect 78932 380156 78988 380196
rect 78932 373072 78988 380100
rect 78932 372596 78988 372624
rect 79044 379596 79100 379618
rect 79044 373072 79100 379540
rect 79044 372596 79100 372624
rect 79156 379148 79212 379188
rect 79156 373072 79212 379092
rect 79156 372596 79212 372624
rect 79268 378700 79324 378740
rect 79268 373072 79324 378644
rect 79268 372596 79324 372624
rect 79380 378252 79436 378292
rect 79380 373072 79436 378196
rect 79380 372596 79436 372624
rect 79492 377804 79548 377844
rect 79492 373072 79548 377748
rect 79492 372596 79548 372624
rect 79604 377356 79660 377396
rect 79604 373072 79660 377300
rect 79604 372596 79660 372624
rect 79716 376908 79772 376948
rect 79716 373072 79772 376852
rect 79716 372596 79772 372624
rect 79828 376460 79884 376500
rect 79828 373072 79884 376404
rect 79828 372596 79884 372624
rect 79940 376012 79996 376052
rect 79940 373072 79996 375956
rect 79940 372596 79996 372624
rect 80052 373072 80108 381108
rect 82628 381052 82684 381092
rect 80052 372596 80108 372624
rect 80164 380604 80220 380644
rect 80164 373072 80220 380548
rect 82516 380492 82572 380532
rect 80164 372596 80220 372624
rect 80276 380044 80332 380084
rect 80276 373072 80332 379988
rect 82404 379932 82460 379972
rect 80276 372596 80332 372624
rect 80388 379484 80444 379524
rect 80388 373072 80444 379428
rect 82292 379372 82348 379412
rect 80388 372596 80444 372624
rect 80500 379036 80556 379076
rect 80500 373072 80556 378980
rect 82180 378924 82236 378964
rect 80500 372596 80556 372624
rect 80612 378588 80668 378628
rect 80612 373072 80668 378532
rect 82068 378476 82124 378516
rect 80612 372596 80668 372624
rect 80724 378140 80780 378180
rect 80724 373072 80780 378084
rect 81956 378028 82012 378068
rect 80724 372596 80780 372624
rect 80836 377692 80892 377732
rect 80836 373072 80892 377636
rect 81844 377580 81900 377620
rect 80836 372596 80892 372624
rect 80948 377244 81004 377284
rect 80948 373072 81004 377188
rect 81732 377132 81788 377172
rect 80948 372596 81004 372624
rect 81060 376796 81116 376836
rect 81060 373072 81116 376740
rect 81620 376684 81676 376724
rect 81060 372596 81116 372624
rect 81172 376348 81228 376388
rect 81172 373072 81228 376292
rect 81508 376236 81564 376276
rect 81172 372596 81228 372624
rect 81284 375900 81340 375940
rect 81284 373072 81340 375844
rect 81284 372596 81340 372624
rect 81396 375788 81452 375828
rect 81396 373072 81452 375732
rect 81396 372596 81452 372624
rect 81508 373072 81564 376180
rect 81508 372596 81564 372624
rect 81620 373072 81676 376628
rect 81620 372596 81676 372624
rect 81732 373072 81788 377076
rect 81732 372596 81788 372624
rect 81844 373072 81900 377524
rect 81844 372596 81900 372624
rect 81956 373072 82012 377972
rect 81956 372596 82012 372624
rect 82068 373072 82124 378420
rect 82068 372596 82124 372624
rect 82180 373072 82236 378868
rect 82180 372596 82236 372624
rect 82292 373072 82348 379316
rect 82292 372596 82348 372624
rect 82404 373072 82460 379876
rect 82404 372596 82460 372624
rect 82516 373072 82572 380436
rect 82516 372596 82572 372624
rect 82628 373072 82684 380996
rect 82628 372596 82684 372624
rect 82740 380940 82796 380980
rect 82740 373072 82796 380884
rect 85428 380828 85484 380868
rect 82740 372596 82796 372624
rect 82852 380380 82908 380420
rect 82852 373072 82908 380324
rect 82852 372596 82908 372624
rect 82964 379820 83020 379860
rect 82964 373072 83020 379764
rect 82964 372596 83020 372624
rect 83076 379260 83132 379300
rect 83076 373072 83132 379204
rect 83076 372596 83132 372624
rect 83188 378812 83244 378852
rect 83188 373072 83244 378756
rect 83188 372596 83244 372624
rect 83300 378364 83356 378404
rect 83300 373072 83356 378308
rect 83300 372596 83356 372624
rect 83412 377916 83468 377956
rect 83412 373072 83468 377860
rect 83412 372596 83468 372624
rect 83524 377468 83580 377508
rect 83524 373072 83580 377412
rect 83524 372596 83580 372624
rect 83636 377020 83692 377060
rect 83636 373072 83692 376964
rect 83636 372596 83692 372624
rect 83748 376572 83804 376612
rect 83748 373072 83804 376516
rect 83748 372596 83804 372624
rect 83860 376124 83916 376164
rect 83860 373072 83916 376068
rect 83860 372596 83916 372624
rect 83972 375676 84028 375716
rect 83972 373072 84028 375620
rect 83972 372596 84028 372624
rect 85428 373072 85484 380772
rect 332100 380778 332806 380830
rect 85428 372596 85484 372624
rect 85652 380268 85708 380308
rect 85652 373072 85708 380212
rect 332100 380250 332154 380778
rect 332744 380250 332806 380778
rect 332100 380188 332806 380250
rect 85652 372596 85708 372624
rect 85876 379708 85932 379748
rect 85876 373072 85932 379652
rect 427200 375800 442000 376000
rect 427200 374200 427400 375800
rect 441800 374200 442000 375800
rect 427200 374000 442000 374200
rect 444000 375800 458800 376000
rect 444000 374200 444200 375800
rect 458600 374200 458800 375800
rect 444000 374000 458800 374200
rect 466800 375800 481600 376000
rect 466800 374200 467000 375800
rect 481400 374200 481600 375800
rect 466800 374000 481600 374200
rect 470200 373500 470900 373600
rect 470200 373000 470300 373500
rect 470800 373000 470900 373500
rect 470200 372900 470900 373000
rect 471400 373500 472100 373600
rect 471400 373000 471500 373500
rect 472000 373000 472100 373500
rect 471400 372900 472100 373000
rect 85876 372596 85932 372624
rect 88381 371234 88424 371290
rect 88480 371234 331600 371290
rect 87084 370982 87164 371038
rect 87220 370982 331348 371038
rect 68924 370730 68964 370786
rect 69020 370730 199304 370786
rect 199360 370730 199400 370786
rect 68812 370486 68852 370542
rect 68908 370486 206864 370542
rect 206920 370486 206960 370542
rect 88636 370242 88676 370298
rect 88732 370242 209258 370298
rect 209314 370242 209354 370298
rect 88888 369998 88928 370054
rect 88984 369998 229796 370054
rect 229852 369998 229892 370054
rect 89140 369754 89180 369810
rect 89236 369754 230048 369810
rect 230104 369754 230144 369810
rect 89392 369510 89432 369566
rect 89488 369510 232694 369566
rect 232750 369510 232790 369566
rect 69036 369266 69076 369322
rect 69132 369266 232946 369322
rect 233002 369266 233042 369322
rect 69148 369022 69188 369078
rect 69244 369022 233198 369078
rect 233254 369022 233294 369078
rect 86116 368778 86156 368834
rect 86212 368778 241514 368834
rect 241570 368778 241610 368834
rect 86494 368534 86534 368590
rect 86590 368534 266966 368590
rect 267022 368534 267062 368590
rect 86746 368290 86786 368346
rect 86842 368290 268352 368346
rect 268408 368290 268448 368346
rect 86998 368046 87038 368102
rect 87094 368046 268604 368102
rect 268660 368046 268700 368102
rect 87250 367802 87290 367858
rect 87346 367802 268856 367858
rect 268912 367802 268952 367858
rect 63378 367542 64890 367668
rect 87502 367558 87542 367614
rect 87598 367558 269108 367614
rect 269164 367558 269204 367614
rect 63378 366912 63504 367542
rect 64764 366912 64890 367542
rect 87754 367314 87794 367370
rect 87850 367314 269360 367370
rect 269416 367314 269456 367370
rect 88006 367070 88046 367126
rect 88102 367070 269612 367126
rect 269668 367070 269708 367126
rect 63378 366786 64890 366912
rect 88258 366826 88298 366882
rect 88354 366826 269864 366882
rect 269920 366826 269960 366882
rect 88510 366582 88550 366638
rect 88606 366582 270116 366638
rect 270172 366582 270212 366638
rect 88762 366338 88802 366394
rect 88858 366338 270368 366394
rect 270424 366338 270464 366394
rect 68252 366094 68292 366150
rect 68348 366094 84980 366150
rect 85036 366094 88480 366150
rect 89014 366094 89054 366150
rect 89110 366094 270620 366150
rect 270676 366094 270716 366150
rect 33400 365800 34800 366000
rect 88424 365906 88480 366094
rect 88424 365850 268100 365906
rect 268156 365850 268179 365906
rect 270832 365850 270872 365906
rect 270928 365850 276220 365906
rect 68476 365606 68516 365662
rect 68572 365606 271124 365662
rect 271180 365606 271220 365662
rect 69260 365362 69300 365418
rect 69356 365362 271376 365418
rect 271432 365362 271472 365418
rect 90428 365118 90468 365174
rect 90524 365118 271628 365174
rect 271684 365118 271724 365174
rect 69616 364874 69636 364930
rect 69692 364874 271880 364930
rect 271936 364874 271976 364930
rect 69508 364630 69524 364686
rect 69580 364630 272132 364686
rect 272188 364630 272228 364686
rect 68700 364386 68740 364442
rect 68796 364386 272384 364442
rect 272440 364386 272480 364442
rect 74425 364142 74452 364198
rect 74508 364142 272636 364198
rect 272692 364142 272732 364198
rect 71612 363898 71652 363954
rect 71708 363898 272888 363954
rect 272944 363898 272984 363954
rect 33400 363600 34800 363800
rect 71500 363654 71540 363710
rect 71596 363654 273140 363710
rect 273196 363654 273236 363710
rect 33400 349200 33600 363600
rect 34600 349200 34800 363600
rect 71388 363410 71428 363466
rect 71484 363410 273392 363466
rect 273448 363410 273488 363466
rect 73180 363166 73220 363222
rect 73276 363166 273644 363222
rect 273700 363166 273740 363222
rect 73068 362922 73108 362978
rect 73164 362922 273896 362978
rect 273952 362922 273992 362978
rect 72956 362678 72996 362734
rect 73052 362678 274148 362734
rect 274204 362678 274244 362734
rect 276164 362724 276220 365850
rect 320670 365486 322812 365612
rect 320670 364604 320796 365486
rect 322686 364604 322812 365486
rect 328500 365400 329300 365500
rect 328500 364800 328600 365400
rect 329200 364800 329300 365400
rect 328500 364700 329300 364800
rect 320670 364478 322812 364604
rect 328500 364000 329300 364100
rect 291144 363544 319645 363600
rect 319701 363544 319717 363600
rect 291144 362724 291200 363544
rect 328500 363400 328600 364000
rect 329200 363400 329300 364000
rect 276164 362668 291200 362724
rect 291368 363320 320684 363376
rect 320740 363320 320788 363376
rect 291368 362490 291424 363320
rect 328500 363300 329300 363400
rect 69372 362434 69412 362490
rect 69468 362434 274400 362490
rect 274456 362434 274496 362490
rect 274864 362434 274904 362490
rect 274960 362434 291424 362490
rect 291662 362922 319438 362978
rect 68028 362190 68068 362246
rect 68124 362190 274652 362246
rect 274708 362190 274748 362246
rect 291662 362001 291718 362922
rect 292000 362678 292040 362734
rect 292096 362678 319260 362734
rect 292252 362434 292292 362490
rect 292348 362434 319016 362490
rect 309262 362190 309302 362246
rect 309358 362190 318772 362246
rect 268073 361945 268100 362001
rect 268156 361945 291718 362001
rect 309514 361946 309554 362002
rect 309610 361946 318528 362002
rect 66024 361620 66906 361746
rect 71281 361702 71316 361758
rect 71372 361702 275156 361758
rect 275212 361702 275252 361758
rect 309766 361702 309806 361758
rect 309862 361702 318284 361758
rect 65268 360864 65772 360990
rect 65268 360360 65394 360864
rect 65646 360360 65772 360864
rect 65268 360234 65772 360360
rect 66024 360360 66150 361620
rect 66780 360360 66906 361620
rect 72844 361458 72884 361514
rect 72940 361458 275408 361514
rect 275464 361458 275504 361514
rect 310018 361458 310058 361514
rect 310114 361458 318040 361514
rect 84044 361214 84084 361270
rect 84140 361214 310310 361270
rect 310366 361214 310406 361270
rect 84268 360970 84308 361026
rect 84364 360970 310562 361026
rect 310618 360970 310658 361026
rect 316764 360990 317772 361116
rect 84492 360726 84532 360782
rect 84588 360726 310814 360782
rect 310870 360726 310910 360782
rect 316764 360612 316890 360990
rect 317646 360612 317772 360990
rect 84716 360482 84756 360538
rect 84812 360482 311066 360538
rect 311122 360482 311162 360538
rect 316764 360486 317772 360612
rect 66024 360234 66906 360360
rect 85400 360238 85428 360294
rect 85484 360238 311318 360294
rect 311374 360238 311414 360294
rect 85628 359994 85652 360050
rect 85708 359994 311570 360050
rect 311626 359994 311666 360050
rect 85836 359750 85876 359806
rect 85932 359750 311822 359806
rect 311878 359750 311918 359806
rect 64052 359493 64092 359549
rect 64148 359493 68068 359549
rect 68124 359493 68164 359549
rect 93340 359506 93380 359562
rect 93436 359506 312074 359562
rect 312130 359506 312170 359562
rect 64724 359269 64764 359325
rect 64820 359269 68292 359325
rect 68348 359269 68388 359325
rect 110140 359262 110180 359318
rect 110236 359262 312326 359318
rect 312382 359262 312422 359318
rect 65010 359045 65050 359101
rect 65106 359045 68516 359101
rect 68572 359045 68612 359101
rect 126940 359018 126980 359074
rect 127036 359018 312578 359074
rect 312634 359018 312674 359074
rect 314302 359018 314342 359074
rect 314398 359018 317756 359074
rect 143740 358774 143780 358830
rect 143836 358774 312830 358830
rect 312886 358774 312926 358830
rect 314554 358774 314594 358830
rect 314650 358774 317512 358830
rect 63000 358470 63504 358596
rect 200540 358530 200580 358586
rect 200636 358530 313082 358586
rect 313138 358530 313178 358586
rect 314806 358530 314846 358586
rect 314902 358530 317268 358586
rect 63000 358092 63126 358470
rect 63378 358092 63504 358470
rect 217340 358286 217380 358342
rect 217436 358286 313334 358342
rect 313390 358286 313430 358342
rect 315058 358286 315098 358342
rect 315154 358286 317024 358342
rect 63000 357966 63504 358092
rect 244140 358042 244180 358098
rect 244236 358042 313586 358098
rect 313642 358042 313682 358098
rect 315310 358042 315350 358098
rect 315406 358042 316780 358098
rect 260940 357798 260980 357854
rect 261036 357798 313838 357854
rect 313894 357798 313934 357854
rect 315562 357798 315602 357854
rect 315658 357798 316536 357854
rect 277740 357554 277780 357610
rect 277836 357554 314090 357610
rect 314146 357554 314186 357610
rect 315814 357554 315854 357610
rect 315910 357554 316292 357610
rect 69701 357066 69748 357122
rect 69804 357066 90749 357122
rect 69820 356822 69860 356878
rect 69916 356822 90749 356878
rect 70044 356578 70084 356634
rect 70140 356578 90846 356634
rect 69932 356334 69972 356390
rect 70028 356334 90846 356390
rect 73292 356090 73332 356146
rect 73388 356090 89824 356146
rect 90170 356090 90720 356146
rect 73404 355846 73444 355902
rect 73500 355846 89824 355902
rect 90170 355846 90846 355902
rect 73516 355602 73556 355658
rect 73612 355602 89824 355658
rect 90170 355602 90846 355658
rect 73628 355358 73668 355414
rect 73724 355358 89824 355414
rect 90170 355358 90846 355414
rect 73740 355114 73780 355170
rect 73836 355114 89824 355170
rect 90170 355114 90846 355170
rect 73852 354870 73892 354926
rect 73948 354870 89824 354926
rect 90170 354870 90846 354926
rect 73964 354626 74004 354682
rect 74060 354626 89824 354682
rect 90170 354626 90846 354682
rect 74076 354382 74116 354438
rect 74172 354382 89824 354438
rect 90170 354382 90846 354438
rect 74188 354138 74228 354194
rect 74284 354138 89824 354194
rect 90170 354138 90846 354194
rect 74300 353894 74340 353950
rect 74396 353894 89824 353950
rect 90170 353894 90846 353950
rect 71164 353650 71204 353706
rect 71260 353650 90846 353706
rect 71052 353406 71092 353462
rect 71148 353406 90846 353462
rect 70940 353162 70980 353218
rect 71036 353162 90846 353218
rect 70828 352918 70868 352974
rect 70924 352918 90846 352974
rect 70716 352674 70756 352730
rect 70812 352674 90846 352730
rect 70604 352430 70644 352486
rect 70700 352430 90846 352486
rect 70492 352186 70532 352242
rect 70588 352186 90846 352242
rect 70380 351942 70420 351998
rect 70476 351942 90846 351998
rect 70268 351698 70308 351754
rect 70364 351698 90846 351754
rect 70156 351454 70196 351510
rect 70252 351454 90846 351510
rect 71724 351210 71764 351266
rect 71820 351210 90846 351266
rect 71836 350966 71876 351022
rect 71932 350966 90846 351022
rect 71948 350722 71988 350778
rect 72044 350722 90846 350778
rect 72060 350478 72100 350534
rect 72156 350478 90846 350534
rect 72172 350234 72212 350290
rect 72268 350234 90846 350290
rect 72284 349990 72324 350046
rect 72380 349990 90846 350046
rect 72396 349746 72436 349802
rect 72492 349746 90846 349802
rect 72508 349502 72548 349558
rect 72604 349502 90874 349558
rect 72620 349258 72660 349314
rect 72716 349258 90720 349314
rect 33400 349000 34800 349200
rect 72732 349014 72772 349070
rect 72828 349014 90846 349070
rect 85610 348770 86912 348826
rect 86968 348770 90846 348826
rect 84940 348526 84980 348582
rect 85036 348526 90846 348582
rect 85621 348282 86408 348338
rect 86464 348282 90846 348338
rect 85318 348038 85358 348094
rect 85414 348038 90846 348094
rect 85619 347794 88172 347850
rect 88228 347794 90846 347850
rect 85617 347550 86660 347606
rect 86716 347550 90846 347606
rect 85619 347306 87668 347362
rect 87724 347306 90846 347362
rect 85615 347062 87416 347118
rect 87472 347062 90846 347118
rect 85610 346818 87920 346874
rect 87976 346818 90846 346874
rect 85052 346574 85092 346630
rect 85148 346574 90846 346630
rect 34570 336980 34580 337036
rect 34636 336980 68516 337036
rect 68572 336980 68582 337036
rect 316236 336540 316292 357554
rect 316480 336784 316536 357798
rect 316724 337028 316780 358042
rect 316968 337272 317024 358286
rect 317212 337516 317268 358530
rect 317456 337760 317512 358774
rect 317700 338004 317756 359018
rect 317984 338288 318040 361458
rect 318228 338532 318284 361702
rect 318472 338776 318528 361946
rect 318716 339020 318772 362190
rect 318960 339264 319016 362434
rect 319204 339508 319260 362678
rect 319382 360515 319438 362922
rect 321930 362502 323442 362628
rect 321930 361872 322056 362502
rect 323316 361872 323442 362502
rect 321930 361746 323442 361872
rect 319380 360360 319438 360515
rect 319380 339676 319436 360360
rect 331292 360328 331348 370982
rect 331544 360454 331600 371234
rect 472400 363600 478000 363800
rect 334400 362200 346200 362400
rect 334400 360800 334600 362200
rect 346000 360800 346200 362200
rect 334400 360600 346200 360800
rect 331544 360398 351130 360454
rect 331292 360272 351004 360328
rect 350948 342310 351004 360272
rect 351074 342436 351130 360398
rect 472400 349200 472600 363600
rect 477800 349200 478000 363600
rect 472400 349000 478000 349200
rect 351074 342380 410640 342436
rect 410700 342380 410740 342436
rect 350948 342254 410800 342310
rect 410860 342254 410906 342310
rect 410130 341712 412020 341838
rect 410130 340578 410256 341712
rect 411894 340578 412020 341712
rect 410130 340452 412020 340578
rect 319380 339620 396116 339676
rect 396172 339620 482160 339676
rect 482216 339620 482236 339676
rect 319204 339452 480410 339508
rect 480466 339452 480506 339508
rect 318960 339208 480158 339264
rect 480214 339208 480254 339264
rect 318716 338964 479906 339020
rect 479962 338964 480002 339020
rect 318472 338720 479654 338776
rect 479710 338720 479750 338776
rect 318228 338476 479402 338532
rect 479458 338476 479498 338532
rect 317984 338232 479150 338288
rect 479206 338232 479246 338288
rect 317700 337948 478898 338004
rect 478954 337948 478994 338004
rect 317456 337704 478646 337760
rect 478702 337704 478742 337760
rect 317212 337460 480662 337516
rect 480718 337460 480758 337516
rect 316968 337216 481670 337272
rect 481726 337216 481766 337272
rect 316724 336972 481418 337028
rect 481474 336972 481514 337028
rect 316480 336728 481166 336784
rect 481222 336728 481262 336784
rect 316236 336484 480914 336540
rect 480970 336484 481010 336540
rect 33078 336226 33506 336260
rect 33078 335888 33120 336226
rect 33462 335888 33506 336226
rect 316134 336204 465290 336260
rect 465346 336204 465386 336260
rect 316106 335960 461510 336016
rect 461566 335960 461606 336016
rect 33078 335846 33506 335888
rect 316134 335716 457730 335772
rect 457786 335716 457866 335772
rect 316134 335472 454076 335528
rect 454132 335472 454172 335528
rect 316134 335228 450296 335284
rect 450352 335228 450392 335284
rect 316106 334984 446516 335040
rect 446572 334984 446612 335040
rect 316134 334740 442736 334796
rect 442792 334740 442832 334796
rect 316134 334496 438956 334552
rect 439012 334496 439052 334552
rect 316134 334252 435176 334308
rect 435232 334252 435272 334308
rect 316134 334008 431396 334064
rect 431452 334008 431492 334064
rect 316134 333764 427616 333820
rect 427672 333764 427712 333820
rect 316134 333520 423962 333576
rect 424018 333520 424058 333576
rect 316134 333276 420182 333332
rect 420238 333276 420278 333332
rect 316106 333032 416402 333088
rect 416458 333032 416498 333088
rect 316134 332788 412622 332844
rect 412678 332788 412718 332844
rect 316134 332544 408842 332600
rect 408898 332544 408938 332600
rect 316134 332300 389438 332356
rect 389494 332300 389534 332356
rect 316106 332056 385658 332112
rect 385714 332056 385754 332112
rect 316134 331812 381878 331868
rect 381934 331812 381974 331868
rect 316134 331568 378098 331624
rect 378154 331568 378194 331624
rect 316134 331324 374318 331380
rect 374374 331324 374414 331380
rect 316134 331080 370538 331136
rect 370594 331080 370634 331136
rect 316134 330836 366758 330892
rect 366814 330836 366854 330892
rect 316134 330592 363104 330648
rect 363160 330592 363200 330648
rect 316134 330348 359324 330404
rect 359380 330348 359420 330404
rect 316134 330104 355544 330160
rect 355600 330104 355640 330160
rect 316134 329860 351764 329916
rect 351820 329860 351860 329916
rect 316134 329616 347984 329672
rect 348040 329616 351099 329672
rect 316134 329372 344204 329428
rect 344260 329372 349307 329428
rect 316134 329128 340424 329184
rect 340480 329128 350683 329184
rect 316134 328884 336644 328940
rect 336700 328884 336740 328940
rect 316134 328640 332990 328696
rect 333046 328640 339931 328696
rect 316134 328396 439460 328452
rect 439516 328396 443240 328452
rect 443296 328396 447020 328452
rect 447076 328396 450800 328452
rect 450856 328396 454580 328452
rect 454636 328396 458234 328452
rect 458290 328396 462014 328452
rect 462070 328396 465794 328452
rect 465850 328396 465890 328452
rect 316134 328152 409346 328208
rect 409402 328152 413126 328208
rect 413182 328152 416906 328208
rect 416962 328152 420686 328208
rect 420742 328152 424466 328208
rect 424522 328152 428120 328208
rect 428176 328152 431900 328208
rect 431956 328152 435680 328208
rect 435736 328152 435776 328208
rect 316134 327908 363608 327964
rect 363664 327908 367262 327964
rect 367318 327908 371042 327964
rect 371098 327908 374822 327964
rect 374878 327908 378602 327964
rect 378658 327908 382382 327964
rect 382438 327908 386162 327964
rect 386218 327908 389942 327964
rect 389998 327908 390038 327964
rect 316134 327664 333368 327720
rect 333424 327664 337148 327720
rect 337204 327664 340928 327720
rect 340984 327664 344708 327720
rect 344764 327664 348488 327720
rect 348544 327664 352268 327720
rect 352324 327664 356048 327720
rect 356104 327664 359828 327720
rect 359884 327664 379587 327720
rect 316134 327420 404558 327476
rect 404614 327420 404654 327476
rect 316134 327176 404054 327232
rect 404110 327176 404150 327232
rect 316134 326932 401534 326988
rect 401590 326932 401630 326988
rect 316134 326688 396872 326744
rect 396928 326688 396968 326744
rect 316106 326444 398006 326500
rect 398062 326444 398102 326500
rect 316134 326200 402542 326256
rect 402598 326200 402638 326256
rect 316134 325956 402038 326012
rect 402094 325956 402134 326012
rect 316134 325712 403046 325768
rect 403102 325712 403142 325768
rect 316134 325468 403550 325524
rect 403606 325468 403646 325524
rect 316134 325224 405062 325280
rect 405118 325224 405158 325280
rect 316134 324980 405566 325036
rect 405622 324980 405662 325036
rect 316134 324736 406070 324792
rect 406126 324736 406166 324792
rect 316134 324492 333872 324548
rect 333928 324492 378347 324548
rect 316106 324248 337652 324304
rect 337708 324248 337748 324304
rect 316134 324004 341432 324060
rect 341488 324004 341528 324060
rect 316134 323760 345212 323816
rect 345268 323760 378995 323816
rect 316134 323516 348992 323572
rect 349048 323516 349088 323572
rect 316134 323272 352772 323328
rect 352828 323272 352868 323328
rect 316106 323028 356552 323084
rect 356608 323028 356648 323084
rect 316134 322784 360332 322840
rect 360388 322784 360428 322840
rect 316134 322540 364112 322596
rect 364168 322540 364208 322596
rect 316134 322296 367766 322352
rect 367822 322296 376651 322352
rect 316134 322052 371546 322108
rect 371602 322052 371642 322108
rect 316134 321808 375326 321864
rect 375382 321808 375803 321864
rect 316134 321564 379106 321620
rect 379162 321564 379202 321620
rect 316134 321320 382886 321376
rect 382942 321320 382982 321376
rect 316134 321076 386666 321132
rect 386722 321076 386762 321132
rect 316134 320832 390446 320888
rect 390502 320832 390542 320888
rect 316134 320588 409850 320644
rect 409906 320588 409946 320644
rect 316134 320344 413630 320400
rect 413686 320344 413726 320400
rect 316134 320100 417410 320156
rect 417466 320100 417506 320156
rect 316134 319856 421190 319912
rect 421246 319856 421286 319912
rect 316134 319612 424970 319668
rect 425026 319612 425066 319668
rect 316134 319368 428624 319424
rect 428680 319368 428720 319424
rect 316134 319124 432404 319180
rect 432460 319124 432500 319180
rect 316134 318880 436184 318936
rect 436240 318880 436280 318936
rect 316134 318636 439964 318692
rect 440020 318636 440060 318692
rect 316106 318392 443744 318448
rect 443800 318392 443840 318448
rect 316134 318148 447524 318204
rect 447580 318148 447620 318204
rect 316134 317904 451304 317960
rect 451360 317904 451400 317960
rect 85590 317782 86282 317838
rect 86338 317782 90720 317838
rect 316134 317660 455084 317716
rect 455140 317660 455180 317716
rect 85600 317538 89306 317594
rect 89362 317538 90720 317594
rect 316134 317416 458738 317472
rect 458794 317416 458834 317472
rect 85600 317294 89558 317350
rect 89614 317294 90720 317350
rect 316134 317172 462518 317228
rect 462574 317172 462614 317228
rect 85600 317050 89810 317106
rect 89866 317050 90720 317106
rect 316134 316928 466298 316984
rect 466354 316928 466394 316984
rect 85600 316806 89936 316862
rect 89992 316806 90720 316862
rect 316358 316798 316414 316821
rect 85990 316562 86030 316618
rect 86086 316562 90720 316618
rect 316414 316684 395558 316740
rect 395714 316684 395752 316740
rect 316358 316597 316414 316615
rect 85738 316318 85778 316374
rect 85834 316318 90720 316374
rect 85486 316074 85526 316130
rect 85582 316074 90749 316130
rect 85234 315830 85274 315886
rect 85330 315830 90720 315886
rect 84982 315586 85022 315642
rect 85078 315586 90720 315642
rect 84730 315342 84770 315398
rect 84826 315342 90720 315398
rect 84478 315098 84518 315154
rect 84574 315098 90720 315154
rect 36708 315029 36726 315085
rect 36786 315029 44138 315085
rect 44198 315084 62496 315085
rect 44198 315029 62343 315084
rect 62333 315027 62343 315029
rect 62400 315029 62496 315084
rect 62400 315027 62410 315029
rect 65734 314979 65750 315035
rect 65826 314979 66048 315035
rect 66108 314979 66228 315035
rect 66288 314979 66306 315035
rect 41132 314906 41151 314966
rect 41211 314906 46265 314966
rect 46325 314906 46339 314966
rect 48444 314841 68852 314861
rect 42289 314785 42308 314841
rect 42364 314805 68852 314841
rect 68908 314805 68948 314861
rect 84226 314854 84266 314910
rect 84322 314854 90720 314910
rect 42364 314785 48516 314805
rect 41310 314673 41326 314729
rect 41386 314673 46871 314729
rect 46931 314673 47959 314729
rect 48019 314673 48042 314729
rect 48444 314617 68964 314637
rect 42519 314561 42532 314617
rect 42588 314581 68964 314617
rect 69020 314581 69060 314637
rect 85565 314610 85904 314666
rect 85960 314610 90720 314666
rect 42588 314561 48514 314581
rect 49324 314357 49364 314413
rect 49420 314357 69076 314413
rect 69132 314357 69172 314413
rect 85612 314366 85652 314422
rect 85708 314366 90720 314422
rect 49548 314133 49588 314189
rect 49644 314133 69188 314189
rect 69244 314133 69284 314189
rect 85360 314122 85400 314178
rect 85456 314122 90720 314178
rect 36476 313906 36486 313966
rect 36546 313964 38110 313966
rect 64095 313964 69300 313965
rect 36546 313908 62692 313964
rect 62748 313908 62776 313964
rect 64095 313909 64135 313964
rect 36546 313906 38110 313908
rect 64125 313907 64135 313909
rect 64192 313909 69300 313964
rect 69356 313909 69396 313965
rect 64192 313907 64202 313909
rect 85108 313878 85148 313934
rect 85204 313878 90720 313934
rect 35028 313488 36036 313614
rect 35028 312984 35154 313488
rect 35910 312984 36036 313488
rect 38386 313604 38625 313632
rect 38386 313329 38413 313604
rect 38578 313329 38625 313604
rect 39853 313597 40093 313653
rect 39853 313333 39889 313597
rect 40051 313333 40093 313597
rect 41725 313623 41985 313646
rect 41725 313357 41744 313623
rect 41962 313357 41985 313623
rect 41725 313338 41985 313357
rect 42714 313614 43344 313740
rect 35028 312858 36036 312984
rect 39853 312396 40093 313333
rect 42714 312858 42840 313614
rect 43218 312858 43344 313614
rect 43974 313687 44478 313740
rect 43974 313428 44030 313687
rect 44407 313428 44478 313687
rect 63044 313685 63084 313741
rect 63140 313685 69412 313741
rect 69468 313685 69510 313741
rect 43974 313362 44478 313428
rect 45447 313601 45647 313624
rect 45447 313339 45467 313601
rect 45631 313339 45647 313601
rect 45447 313322 45647 313339
rect 46908 313610 47148 313656
rect 46908 313336 46935 313610
rect 47111 313336 47148 313610
rect 48764 313634 49026 313649
rect 84856 313634 84896 313690
rect 84952 313634 90720 313690
rect 48764 313364 48779 313634
rect 49011 313364 49026 313634
rect 48764 313345 49026 313364
rect 60228 313362 61362 313488
rect 65899 313461 65927 313517
rect 65984 313461 69524 313517
rect 69580 313461 69590 313517
rect 84604 313390 84644 313446
rect 84700 313390 90720 313446
rect 42714 312732 43344 312858
rect 46908 312396 47148 313336
rect 60228 313110 60354 313362
rect 61236 313110 61362 313362
rect 67679 313237 67719 313293
rect 67776 313237 69636 313293
rect 69692 313237 69702 313293
rect 84352 313146 84392 313202
rect 84448 313146 90720 313202
rect 60228 312984 61362 313110
rect 64386 312732 65520 312858
rect 64386 312480 64512 312732
rect 65394 312480 65520 312732
rect 39853 312393 50898 312396
rect 39853 312160 50283 312393
rect 50882 312160 50898 312393
rect 64386 312354 65520 312480
rect 39853 312156 50898 312160
rect 56634 312117 56644 312173
rect 56700 312117 68740 312173
rect 68796 312117 68836 312173
rect 60228 311724 61362 311850
rect 60228 311472 60354 311724
rect 61236 311472 61362 311724
rect 60228 311346 61362 311472
rect 68544 311220 69552 311346
rect 68544 310968 68670 311220
rect 69426 310968 69552 311220
rect 42714 310842 43344 310968
rect 42714 310338 42840 310842
rect 43218 310338 43344 310842
rect 42714 310212 43344 310338
rect 49896 310842 50526 310968
rect 68544 310842 69552 310968
rect 49896 310338 50022 310842
rect 50400 310338 50526 310842
rect 64134 310716 64184 310842
rect 64240 310716 64386 310842
rect 65520 310716 65976 310842
rect 66032 310716 67768 310842
rect 67824 310716 67914 310842
rect 64498 310535 64520 310611
rect 64596 310535 67446 310611
rect 67522 310535 67558 310611
rect 49896 310212 50526 310338
rect 57886 310424 58126 310447
rect 57886 310206 57903 310424
rect 58105 310206 58126 310424
rect 57886 310183 58126 310206
rect 50526 309582 51408 309708
rect 50526 309078 50652 309582
rect 51282 309078 51408 309582
rect 50526 308952 51408 309078
rect 58464 309582 58968 309708
rect 58464 308952 58590 309582
rect 58842 308952 58968 309582
rect 58464 308826 58968 308952
rect 32478 308528 32550 308767
rect 32810 308528 38386 308767
rect 38625 308528 45418 308767
rect 45657 308528 52708 308767
rect 52947 308528 52979 308767
rect 33109 308123 33150 308296
rect 33410 308285 51981 308296
rect 33410 308134 51619 308285
rect 51968 308134 51981 308285
rect 33410 308123 51981 308134
rect 84100 305582 84140 305638
rect 84196 305582 90972 305638
rect 32748 286356 32788 286412
rect 32844 286356 82740 286412
rect 82796 286356 82836 286412
rect 33308 286244 33348 286300
rect 33404 286244 82964 286300
rect 83020 286244 83060 286300
rect 33868 286132 33908 286188
rect 33964 286132 83188 286188
rect 83244 286132 83284 286188
rect 34428 286020 34468 286076
rect 34524 286020 83412 286076
rect 83468 286020 83508 286076
rect 34316 285908 34356 285964
rect 34412 285908 76356 285964
rect 76412 285908 76452 285964
rect 33756 285796 33796 285852
rect 33852 285796 76244 285852
rect 76300 285796 76340 285852
rect 33196 285684 33236 285740
rect 33292 285684 76132 285740
rect 76188 285684 76228 285740
rect 32636 285572 32676 285628
rect 32732 285572 76020 285628
rect 76076 285572 76116 285628
rect 34204 285460 34244 285516
rect 34300 285460 75908 285516
rect 75964 285460 76004 285516
rect 33644 285348 33684 285404
rect 33740 285348 75796 285404
rect 75852 285348 75892 285404
rect 33084 285236 33124 285292
rect 33180 285236 75684 285292
rect 75740 285236 75780 285292
rect 32524 285124 32564 285180
rect 32620 285124 75572 285180
rect 75628 285124 75668 285180
rect 34092 285012 34132 285068
rect 34188 285012 75460 285068
rect 75516 285012 75556 285068
rect 33532 284900 33572 284956
rect 33628 284900 75348 284956
rect 75404 284900 75444 284956
rect 32972 284788 33012 284844
rect 33068 284788 75236 284844
rect 75292 284788 75332 284844
rect 32412 284676 32452 284732
rect 32508 284676 75124 284732
rect 75180 284676 75220 284732
rect 33980 284564 34020 284620
rect 34076 284564 75012 284620
rect 75068 284564 75108 284620
rect 33420 284452 33460 284508
rect 33516 284452 74900 284508
rect 74956 284452 74996 284508
rect 32860 284340 32900 284396
rect 32956 284340 74788 284396
rect 74844 284340 74884 284396
rect 32300 284228 32340 284284
rect 32396 284228 74676 284284
rect 74732 284228 74772 284284
rect 48462 283951 50274 284004
rect 48462 283874 49186 283951
rect 33490 283714 33526 283874
rect 33670 283714 49186 283874
rect 48462 283673 49186 283714
rect 50234 283673 50274 283951
rect 48462 283626 50274 283673
rect 54810 283944 56740 284004
rect 54810 283680 54858 283944
rect 55884 283680 56740 283944
rect 54810 283626 56740 283680
rect 48462 283374 49062 283626
rect 56140 283374 56740 283626
rect 56860 283922 68976 284032
rect 69088 283922 69128 284032
rect 56860 283447 57180 283922
rect 34870 281649 34950 282082
rect 35210 282078 38339 282082
rect 35210 281653 37740 282078
rect 38303 281653 38339 282078
rect 35210 281649 38339 281653
rect 82588 266582 82628 266638
rect 82684 266582 90880 266638
rect 82476 260564 82516 260620
rect 82572 260564 90748 260620
rect 82364 260320 82404 260376
rect 82460 260320 90749 260376
rect 82252 260076 82292 260132
rect 82348 260076 90749 260132
rect 82140 259832 82180 259888
rect 82236 259832 90846 259888
rect 82028 259588 82068 259644
rect 82124 259588 90720 259644
rect 81916 259344 81956 259400
rect 82012 259344 90720 259400
rect 81804 259100 81844 259156
rect 81900 259100 90846 259156
rect 81692 258856 81732 258912
rect 81788 258856 90846 258912
rect 81580 258612 81620 258668
rect 81676 258612 90846 258668
rect 81468 258368 81508 258424
rect 81564 258368 90846 258424
rect 81356 258124 81396 258180
rect 81452 258124 90846 258180
rect 76316 257880 76356 257936
rect 76412 257880 90846 257936
rect 76204 257636 76244 257692
rect 76300 257636 90720 257692
rect 76092 257392 76132 257448
rect 76188 257392 90720 257448
rect 33695 257206 34047 257276
rect 33695 254062 33739 257206
rect 33994 254062 34047 257206
rect 75980 257148 76020 257204
rect 76076 257148 90720 257204
rect 75532 256904 75572 256960
rect 75628 256904 90720 256960
rect 75644 256660 75684 256716
rect 75740 256660 90846 256716
rect 75756 256416 75796 256472
rect 75852 256416 90846 256472
rect 75868 256172 75908 256228
rect 75964 256172 90846 256228
rect 81244 255928 81284 255984
rect 81340 255928 90846 255984
rect 81132 255684 81172 255740
rect 81228 255684 90846 255740
rect 81020 255440 81060 255496
rect 81116 255440 90720 255496
rect 80908 255196 80948 255252
rect 81004 255196 90720 255252
rect 80796 254952 80836 255008
rect 80892 254952 90720 255008
rect 80684 254708 80724 254764
rect 80780 254708 90720 254764
rect 80572 254464 80612 254520
rect 80668 254464 90720 254520
rect 80460 254220 80500 254276
rect 80556 254220 90720 254276
rect 33695 254010 34047 254062
rect 80348 253976 80388 254032
rect 80444 253976 90720 254032
rect 80236 253732 80276 253788
rect 80332 253732 90846 253788
rect 80124 253488 80164 253544
rect 80220 253488 90846 253544
rect 80012 253244 80052 253300
rect 80108 253244 90846 253300
rect 79900 253000 79940 253056
rect 79996 253000 90846 253056
rect 79788 252756 79828 252812
rect 79884 252756 90846 252812
rect 79676 252512 79716 252568
rect 79772 252512 90846 252568
rect 79564 252268 79604 252324
rect 79660 252268 90846 252324
rect 79452 252024 79492 252080
rect 79548 252024 90846 252080
rect 79340 251780 79380 251836
rect 79436 251780 90846 251836
rect 79228 251536 79268 251592
rect 79324 251536 90846 251592
rect 79116 251292 79156 251348
rect 79212 251292 90846 251348
rect 79004 251048 79044 251104
rect 79100 251048 90846 251104
rect 78892 250804 78932 250860
rect 78988 250804 90846 250860
rect 78780 250560 78820 250616
rect 78876 250560 90846 250616
rect 78668 250316 78708 250372
rect 78764 250316 90720 250372
rect 75420 250072 75460 250128
rect 75516 250072 90720 250128
rect 75308 249828 75348 249884
rect 75404 249828 90720 249884
rect 75196 249584 75236 249640
rect 75292 249584 90846 249640
rect 35507 248888 35550 249475
rect 35810 249473 38189 249475
rect 35810 248893 37590 249473
rect 38138 248893 38189 249473
rect 75084 249340 75124 249396
rect 75180 249340 90846 249396
rect 78556 249096 78596 249152
rect 78652 249096 90846 249152
rect 35810 248888 38189 248893
rect 78444 248852 78484 248908
rect 78540 248852 90846 248908
rect 78332 248608 78372 248664
rect 78428 248608 90846 248664
rect 78220 248364 78260 248420
rect 78316 248364 90846 248420
rect 78108 248120 78148 248176
rect 78204 248120 90846 248176
rect 58464 247968 59346 248094
rect 58464 247086 58590 247968
rect 59220 247086 59346 247968
rect 77996 247876 78036 247932
rect 78092 247876 90846 247932
rect 77884 247632 77924 247688
rect 77980 247632 90846 247688
rect 77772 247388 77812 247444
rect 77868 247388 90846 247444
rect 77660 247144 77700 247200
rect 77756 247144 90720 247200
rect 58464 246960 59346 247086
rect 77548 246900 77588 246956
rect 77644 246900 90846 246956
rect 77436 246656 77476 246712
rect 77532 246656 90846 246712
rect 60102 246330 60982 246456
rect 77324 246412 77364 246468
rect 77420 246412 90846 246468
rect 60102 245448 60228 246330
rect 60858 245448 60982 246330
rect 74972 246168 75012 246224
rect 75068 246168 90846 246224
rect 74860 245924 74900 245980
rect 74956 245924 90720 245980
rect 74748 245680 74788 245736
rect 74844 245680 90846 245736
rect 60102 245322 60982 245448
rect 74636 245436 74676 245492
rect 74732 245436 90846 245492
rect 54050 243784 54106 244936
rect 46076 243728 46116 243784
rect 46172 243728 54106 243784
rect 54172 243662 54228 244936
rect 47868 243606 47908 243662
rect 47964 243606 54228 243662
rect 54294 243540 54350 244936
rect 49660 243484 49700 243540
rect 49756 243484 54350 243540
rect 54416 243418 54472 244936
rect 51452 243362 51492 243418
rect 51548 243362 54472 243418
rect 54538 243296 54594 244936
rect 53244 243240 53284 243296
rect 53340 243240 54594 243296
rect 54660 243174 54716 244936
rect 54782 243296 54838 244936
rect 54904 243418 54960 244936
rect 55026 243540 55082 244936
rect 55148 243662 55204 244936
rect 55270 243784 55326 244936
rect 63756 244692 64764 244818
rect 63756 243936 63882 244692
rect 64638 243936 64764 244692
rect 63756 243882 64764 243936
rect 55270 243748 64036 243784
rect 55272 243728 64036 243748
rect 64092 243728 64132 243784
rect 55148 243606 62244 243662
rect 62300 243606 62340 243662
rect 55026 243484 60452 243540
rect 60508 243484 60548 243540
rect 54904 243362 58660 243418
rect 58716 243362 58756 243418
rect 54782 243240 56868 243296
rect 56924 243240 56964 243296
rect 67158 243180 68040 243306
rect 54660 243118 55076 243174
rect 55132 243118 55152 243174
rect 67158 242298 67284 243180
rect 67914 242298 68040 243180
rect 67158 242172 68040 242298
rect 65638 241794 67024 241920
rect 65638 241290 65764 241794
rect 66898 241290 67024 241794
rect 65638 241164 67024 241290
rect 46076 240816 46116 240872
rect 46172 240816 73332 240872
rect 73388 240816 73428 240872
rect 47868 240694 47908 240750
rect 47964 240694 73444 240750
rect 73500 240694 73540 240750
rect 49660 240572 49700 240628
rect 49756 240572 73556 240628
rect 73612 240572 73652 240628
rect 34295 240406 34647 240476
rect 51452 240450 51492 240506
rect 51548 240450 73668 240506
rect 73724 240450 73764 240506
rect 34295 237262 34339 240406
rect 34594 237262 34647 240406
rect 53244 240328 53284 240384
rect 53340 240328 73780 240384
rect 73836 240328 73876 240384
rect 55036 240206 55076 240262
rect 55132 240206 73892 240262
rect 73948 240206 73988 240262
rect 56828 240084 56868 240140
rect 56924 240084 74004 240140
rect 74060 240084 74100 240140
rect 49644 239904 51786 240030
rect 58620 239962 58660 240018
rect 58716 239962 74116 240018
rect 74172 239962 74212 240018
rect 49644 239778 49770 239904
rect 51660 239778 51786 239904
rect 60412 239840 60452 239896
rect 60508 239840 74228 239896
rect 74284 239840 74324 239896
rect 49644 239652 51786 239778
rect 62204 239718 62244 239774
rect 62300 239718 74340 239774
rect 74396 239718 74436 239774
rect 63996 239596 64036 239652
rect 64092 239596 74452 239652
rect 74508 239596 74548 239652
rect 64849 239346 65109 239378
rect 64849 238630 64857 239346
rect 65097 238630 65109 239346
rect 34870 237449 34950 237882
rect 35210 237878 38339 237882
rect 35210 237453 37740 237878
rect 38303 237453 38339 237878
rect 35210 237449 38339 237453
rect 34295 237210 34647 237262
rect 64849 234149 65109 238630
rect 64849 233949 65109 233982
rect 66276 233604 66780 233730
rect 66276 232596 66402 233604
rect 66654 232596 66780 233604
rect 66276 232470 66780 232596
rect 72324 229320 73710 229446
rect 72324 228690 72450 229320
rect 73584 228690 73710 229320
rect 72324 228564 73710 228690
rect 65268 226795 66654 226800
rect 64213 226767 66654 226795
rect 64213 225689 64234 226767
rect 64745 226674 66654 226767
rect 64745 225792 65394 226674
rect 66528 225792 66654 226674
rect 64745 225689 66654 225792
rect 64213 225666 66654 225689
rect 64213 225664 66526 225666
rect 33126 223223 33425 223279
rect 33126 219357 33176 223223
rect 33382 219357 33425 223223
rect 33126 219314 33425 219357
rect 72828 209538 73710 209664
rect 72828 208656 72954 209538
rect 73584 208656 73710 209538
rect 72828 208530 73710 208656
rect 79254 207942 79758 208026
rect 79254 206980 79331 207942
rect 79685 206980 79758 207942
rect 79254 206892 79758 206980
rect 34895 206806 35247 206876
rect 34895 203662 34939 206806
rect 35194 203662 35247 206806
rect 73404 206658 73444 206714
rect 73500 206658 81956 206714
rect 82012 206658 82052 206714
rect 74076 206546 74116 206602
rect 74172 206546 82068 206602
rect 82124 206546 82164 206602
rect 74748 206434 74788 206490
rect 74844 206434 82180 206490
rect 82236 206434 82276 206490
rect 75420 206322 75460 206378
rect 75516 206322 82292 206378
rect 82348 206322 82388 206378
rect 76092 206210 76132 206266
rect 76188 206210 82404 206266
rect 82460 206210 82500 206266
rect 76764 206098 76804 206154
rect 76860 206098 82516 206154
rect 82572 206098 82612 206154
rect 73768 205944 73780 206000
rect 73836 205944 75124 206000
rect 75180 205944 75200 206000
rect 77436 205986 77476 206042
rect 77532 205986 82628 206042
rect 82684 205986 82724 206042
rect 35507 205288 35550 205875
rect 35810 205873 38189 205875
rect 78108 205874 78148 205930
rect 78204 205874 82740 205930
rect 82796 205874 82836 205930
rect 35810 205293 37590 205873
rect 38138 205293 38189 205873
rect 78780 205762 78820 205818
rect 78876 205762 82852 205818
rect 82908 205762 82948 205818
rect 35810 205288 38189 205293
rect 74306 205722 74654 205762
rect 74306 205038 74345 205722
rect 74614 205038 74654 205722
rect 79452 205650 79492 205706
rect 79548 205650 82964 205706
rect 83020 205650 83060 205706
rect 80124 205538 80164 205594
rect 80220 205538 83076 205594
rect 83132 205538 83172 205594
rect 77340 205426 77364 205482
rect 77420 205426 83188 205482
rect 83244 205426 83284 205482
rect 75530 205314 75572 205370
rect 75628 205314 83300 205370
rect 83356 205314 83396 205370
rect 75084 205202 75124 205258
rect 75180 205202 83412 205258
rect 83468 205202 83508 205258
rect 74306 204996 74654 205038
rect 34895 203610 35247 203662
rect 72344 203634 80164 203690
rect 80220 203634 80258 203690
rect 72344 203512 77364 203568
rect 77420 203512 77452 203568
rect 72344 203390 75572 203446
rect 75628 203390 75668 203446
rect 72344 203268 73780 203324
rect 73836 203268 73876 203324
rect 72344 203146 79492 203202
rect 79548 203146 79588 203202
rect 72344 203024 78820 203080
rect 78876 203024 78916 203080
rect 72344 202902 78148 202958
rect 78204 202902 78244 202958
rect 72344 202780 77476 202836
rect 77532 202780 77558 202836
rect 72344 202658 76804 202714
rect 76860 202658 76900 202714
rect 72344 202536 76132 202592
rect 76188 202536 76228 202592
rect 72344 202414 75460 202470
rect 75516 202414 75556 202470
rect 72344 202292 74788 202348
rect 74844 202292 74884 202348
rect 72344 202170 74116 202226
rect 74172 202170 74194 202226
rect 72344 202048 73444 202104
rect 73500 202048 73540 202104
rect 73080 200970 73836 201096
rect 73080 199710 73206 200970
rect 73710 199710 73836 200970
rect 73080 199584 73836 199710
rect 33715 198886 33750 199085
rect 34010 198886 67957 199085
rect 32438 198151 32550 198350
rect 32810 198151 64545 198350
rect 64831 198151 64885 198350
rect 36046 197377 36150 197670
rect 36410 197377 65443 197670
rect 65722 197377 65798 197670
rect 49789 197117 51889 197164
rect 49789 196869 49829 197117
rect 51830 196869 51889 197117
rect 49789 196826 51889 196869
rect 34870 194649 34950 195082
rect 35210 195078 38339 195082
rect 35210 194653 37740 195078
rect 38303 194653 38339 195078
rect 35210 194649 38339 194653
rect 35495 190006 35847 190076
rect 35495 186862 35539 190006
rect 35794 186862 35847 190006
rect 66024 190008 66906 190134
rect 66024 189252 66150 190008
rect 66780 189252 66906 190008
rect 66024 189126 66906 189252
rect 35495 186810 35847 186862
rect 67758 185993 67957 198886
rect 70686 198850 71442 198976
rect 70686 198094 70812 198850
rect 71316 198094 71442 198850
rect 85618 198628 90188 198684
rect 90244 198628 90754 198684
rect 85618 198384 90062 198440
rect 90118 198384 90754 198440
rect 85618 198140 90314 198196
rect 90370 198140 90754 198196
rect 70686 197968 71442 198094
rect 83847 197286 83888 197342
rect 83944 197286 90754 197342
rect 68922 193032 69678 193158
rect 68922 192402 69048 193032
rect 69552 192402 69678 193032
rect 68922 192276 69678 192402
rect 66767 185968 67957 185993
rect 66767 185801 66801 185968
rect 67096 185801 67957 185968
rect 66767 185794 67957 185801
rect 66770 185782 67122 185794
rect 64248 182952 64260 184338
rect 64764 184212 67032 184338
rect 64764 183078 65772 184212
rect 66906 183078 67032 184212
rect 64764 182952 67032 183078
rect 36095 173206 36447 173276
rect 36095 170062 36139 173206
rect 36394 170062 36447 173206
rect 36095 170010 36447 170062
rect 73206 167202 74214 167328
rect 73206 166446 73332 167202
rect 74088 166446 74214 167202
rect 73206 166320 74214 166446
rect 79380 165312 80010 165438
rect 79380 164178 79506 165312
rect 79884 164178 80010 165312
rect 79380 164052 80010 164178
rect 73404 163836 73444 163892
rect 73500 163836 80388 163892
rect 80444 163836 80484 163892
rect 74076 163724 74116 163780
rect 74172 163724 80500 163780
rect 80556 163724 80596 163780
rect 74748 163612 74788 163668
rect 74844 163612 80612 163668
rect 80668 163612 80708 163668
rect 75420 163500 75460 163556
rect 75516 163500 80724 163556
rect 80780 163500 80820 163556
rect 76092 163388 76132 163444
rect 76188 163388 80836 163444
rect 80892 163388 80932 163444
rect 76764 163276 76804 163332
rect 76860 163276 80948 163332
rect 81004 163276 81044 163332
rect 77436 163164 77476 163220
rect 77532 163164 81060 163220
rect 81116 163164 81156 163220
rect 35507 162488 35550 163075
rect 35810 163073 38189 163075
rect 35810 162493 37590 163073
rect 38138 162493 38189 163073
rect 78108 163052 78148 163108
rect 78204 163052 81172 163108
rect 81228 163052 81268 163108
rect 78780 162940 78820 162996
rect 78876 162940 81284 162996
rect 81340 162940 81380 162996
rect 79452 162828 79492 162884
rect 79548 162828 81396 162884
rect 81452 162828 81492 162884
rect 80124 162716 80164 162772
rect 80220 162716 81508 162772
rect 81564 162716 81604 162772
rect 77334 162604 77364 162660
rect 77420 162604 81620 162660
rect 81676 162604 81716 162660
rect 35810 162488 38189 162493
rect 75550 162492 75572 162548
rect 75628 162492 81732 162548
rect 81788 162492 81828 162548
rect 73738 162380 73780 162436
rect 73836 162380 81844 162436
rect 81900 162380 81933 162436
rect 80766 162036 81648 162162
rect 80766 161532 80892 162036
rect 81522 161532 81648 162036
rect 80766 161406 81648 161532
rect 72344 160812 80164 160868
rect 80220 160812 80230 160868
rect 72344 160690 77364 160746
rect 77420 160690 77452 160746
rect 72344 160568 75572 160624
rect 75628 160568 75668 160624
rect 72344 160446 73780 160502
rect 73836 160446 73876 160502
rect 72344 160324 79492 160380
rect 79548 160324 79588 160380
rect 72344 160202 78820 160258
rect 78876 160202 78916 160258
rect 72344 160080 78148 160136
rect 78204 160080 78244 160136
rect 72344 159958 77476 160014
rect 77532 159958 77548 160014
rect 72344 159836 76804 159892
rect 76860 159836 76900 159892
rect 72344 159714 76132 159770
rect 76188 159714 76228 159770
rect 72344 159592 75460 159648
rect 75516 159592 75556 159648
rect 72344 159470 74788 159526
rect 74844 159470 74884 159526
rect 72344 159348 74116 159404
rect 74172 159348 74206 159404
rect 72344 159226 73444 159282
rect 73500 159226 73540 159282
rect 70878 156752 71846 156878
rect 70878 156500 70964 156752
rect 71720 156500 71846 156752
rect 36695 156406 37047 156476
rect 36695 153262 36739 156406
rect 36994 153262 37047 156406
rect 70878 156374 71846 156500
rect 71986 156744 72954 156870
rect 71986 156492 72072 156744
rect 72828 156492 72954 156744
rect 71986 156366 72954 156492
rect 61674 155540 61684 155596
rect 61740 155540 83748 155596
rect 83804 155540 83830 155596
rect 59964 155400 60004 155456
rect 60060 155400 83888 155456
rect 83944 155400 83964 155456
rect 61756 155278 61796 155334
rect 61852 155278 84014 155334
rect 84070 155278 84087 155334
rect 62316 155156 62356 155212
rect 62412 155156 84140 155212
rect 84196 155156 84236 155212
rect 62428 155034 62468 155090
rect 62524 155034 84266 155090
rect 84322 155034 84362 155090
rect 62988 154912 63028 154968
rect 63084 154912 84392 154968
rect 84448 154912 84488 154968
rect 63100 154790 63140 154846
rect 63196 154790 84518 154846
rect 84574 154790 84614 154846
rect 63660 154668 63700 154724
rect 63756 154668 84644 154724
rect 84700 154668 84740 154724
rect 63772 154546 63812 154602
rect 63868 154546 84770 154602
rect 84826 154546 84866 154602
rect 64332 154424 64372 154480
rect 64428 154424 84896 154480
rect 84952 154424 84992 154480
rect 64444 154302 64484 154358
rect 64540 154302 85022 154358
rect 85078 154302 85118 154358
rect 65004 154180 65044 154236
rect 65100 154180 85148 154236
rect 85204 154180 85244 154236
rect 65116 154058 65156 154114
rect 65212 154058 85274 154114
rect 85330 154058 85370 154114
rect 65676 153936 65716 153992
rect 65772 153936 85400 153992
rect 85456 153936 85496 153992
rect 65788 153814 65828 153870
rect 65884 153814 85526 153870
rect 85582 153814 85622 153870
rect 66348 153692 66388 153748
rect 66444 153692 85652 153748
rect 85708 153692 85748 153748
rect 36695 153210 37047 153262
rect 51282 153468 52920 153594
rect 66460 153570 66500 153626
rect 66556 153570 85778 153626
rect 85834 153570 85874 153626
rect 51282 152838 51408 153468
rect 52794 152838 52920 153468
rect 67020 153448 67060 153504
rect 67116 153448 85904 153504
rect 85960 153448 86000 153504
rect 67132 153326 67172 153382
rect 67228 153326 86030 153382
rect 86086 153326 86126 153382
rect 67692 153204 67732 153260
rect 67788 153204 86156 153260
rect 86212 153204 86252 153260
rect 67804 153082 67844 153138
rect 67900 153082 86282 153138
rect 86338 153082 86378 153138
rect 86134 152960 86156 153016
rect 86212 152960 87164 153016
rect 87220 152960 87230 153016
rect 68364 152838 68404 152894
rect 68460 152838 86534 152894
rect 86590 152838 86630 152894
rect 51282 152712 52920 152838
rect 68810 152716 68850 152772
rect 68910 152716 86660 152772
rect 86716 152716 86756 152772
rect 69036 152594 69076 152650
rect 69132 152594 86786 152650
rect 86842 152594 86882 152650
rect 69596 152472 69636 152528
rect 69692 152472 86912 152528
rect 86968 152472 87008 152528
rect 69708 152350 69748 152406
rect 69804 152350 87038 152406
rect 87094 152350 87134 152406
rect 70268 152228 70308 152284
rect 70364 152228 87164 152284
rect 87220 152228 87260 152284
rect 70380 152106 70420 152162
rect 70476 152106 87290 152162
rect 87346 152106 87386 152162
rect 70940 151984 70980 152040
rect 71036 151984 87416 152040
rect 87472 151984 87512 152040
rect 71052 151862 71092 151918
rect 71148 151862 87542 151918
rect 87598 151862 87638 151918
rect 71612 151740 71652 151796
rect 71708 151740 87668 151796
rect 87724 151740 87764 151796
rect 71724 151618 71764 151674
rect 71820 151618 87794 151674
rect 87850 151618 87890 151674
rect 72284 151496 72324 151552
rect 72380 151496 87920 151552
rect 87976 151496 88016 151552
rect 72396 151374 72436 151430
rect 72492 151374 88046 151430
rect 88102 151374 88142 151430
rect 72956 151252 72996 151308
rect 73052 151252 88172 151308
rect 88228 151252 88268 151308
rect 73068 151130 73108 151186
rect 73164 151130 88298 151186
rect 88354 151130 88394 151186
rect 73628 151008 73668 151064
rect 73724 151008 88046 151064
rect 88102 151008 88142 151064
rect 73740 150886 73780 150942
rect 73836 150886 88550 150942
rect 88606 150886 88646 150942
rect 74300 150764 74340 150820
rect 74396 150764 88676 150820
rect 88732 150764 88772 150820
rect 74412 150642 74452 150698
rect 74508 150642 88802 150698
rect 88858 150642 88898 150698
rect 74972 150520 75012 150576
rect 75068 150520 88928 150576
rect 88984 150520 89024 150576
rect 75084 150398 75124 150454
rect 75180 150398 89054 150454
rect 89110 150398 89150 150454
rect 75644 150276 75684 150332
rect 75740 150276 89180 150332
rect 89236 150276 89276 150332
rect 75756 150154 75796 150210
rect 75852 150154 89306 150210
rect 89362 150154 89402 150210
rect 76316 150032 76356 150088
rect 76412 150032 89432 150088
rect 89488 150032 89528 150088
rect 76428 149910 76468 149966
rect 76524 149910 89558 149966
rect 89614 149910 89654 149966
rect 76988 149788 77028 149844
rect 77084 149788 89684 149844
rect 89740 149788 89780 149844
rect 321000 149736 321600 149836
rect 77100 149666 77140 149722
rect 77196 149666 89810 149722
rect 89866 149666 89906 149722
rect 77772 149544 77812 149600
rect 77868 149544 89936 149600
rect 89992 149544 90032 149600
rect 78444 149422 78484 149478
rect 78540 149422 90062 149478
rect 90118 149422 90158 149478
rect 79116 149300 79156 149356
rect 79212 149300 90188 149356
rect 90244 149300 90284 149356
rect 321000 149336 321100 149736
rect 321500 149336 321600 149736
rect 321000 149236 321600 149336
rect 79788 149178 79828 149234
rect 79884 149178 90314 149234
rect 90370 149178 90410 149234
rect 321000 148736 321600 148836
rect 321000 148336 321100 148736
rect 321500 148336 321600 148736
rect 214132 148202 214172 148258
rect 214228 148202 292670 148258
rect 292726 148202 292766 148258
rect 321000 148236 321600 148336
rect 80460 148080 80500 148136
rect 80556 148080 202832 148136
rect 202888 148080 202898 148136
rect 233570 147958 233610 148014
rect 233666 147958 292922 148014
rect 292978 147958 293018 148014
rect 80796 147836 80836 147892
rect 80892 147836 202580 147892
rect 202636 147836 316358 147892
rect 316414 147836 316424 147892
rect 89674 147714 89684 147770
rect 89740 147714 295694 147770
rect 295750 147714 295760 147770
rect 87164 147648 87220 147658
rect 84830 147588 84870 147644
rect 84926 147588 86156 147644
rect 86212 147588 86242 147644
rect 87220 147592 201194 147648
rect 201250 147592 201320 147648
rect 87164 147582 87220 147592
rect 90458 147476 90468 147532
rect 90524 147476 115668 147532
rect 115724 147476 115734 147532
rect 126604 147470 126644 147526
rect 126700 147470 315854 147526
rect 315910 147470 315920 147526
rect 85964 147364 85990 147420
rect 86046 147364 88424 147420
rect 88480 147364 88510 147420
rect 128844 147348 128884 147404
rect 128940 147348 315602 147404
rect 315658 147348 315698 147404
rect 88900 147252 117012 147308
rect 117068 147252 117104 147308
rect 88900 147196 88956 147252
rect 131084 147226 131124 147282
rect 131180 147226 315350 147282
rect 315406 147226 315446 147282
rect 86640 147140 86662 147196
rect 86718 147140 88956 147196
rect 133324 147104 133364 147160
rect 133420 147104 315098 147160
rect 315154 147104 315194 147160
rect 89236 147028 116787 147084
rect 116843 147028 116865 147084
rect 89236 146972 89292 147028
rect 135564 146982 135604 147038
rect 135660 146982 314846 147038
rect 314902 146982 314942 147038
rect 84401 146916 84422 146972
rect 84478 146916 85318 146972
rect 85374 146916 89292 146972
rect 137804 146860 137844 146916
rect 137900 146860 314594 146916
rect 314650 146860 314690 146916
rect 140044 146738 140084 146794
rect 140140 146738 314342 146794
rect 314398 146738 314438 146794
rect 51968 146580 52500 146636
rect 52556 146580 56868 146636
rect 56924 146580 57008 146636
rect 142284 146616 142324 146672
rect 142380 146616 314090 146672
rect 314146 146616 314186 146672
rect 81144 146412 81774 146538
rect 144972 146494 145012 146550
rect 145068 146494 313838 146550
rect 313894 146494 313934 146550
rect 51968 146356 53060 146412
rect 53116 146356 56644 146412
rect 56700 146356 57008 146412
rect 51968 146132 53620 146188
rect 53676 146132 55524 146188
rect 55580 146132 57008 146188
rect 32958 146020 32998 146076
rect 33054 146020 37156 146076
rect 37212 146020 37222 146076
rect 47152 145908 47236 145964
rect 47292 145908 54180 145964
rect 54236 145908 54320 145964
rect 32792 145760 32802 145816
rect 32858 145760 51814 145816
rect 51758 145696 51814 145760
rect 51758 145640 59122 145696
rect 59066 143866 59122 145640
rect 59066 143810 61334 143866
rect 61390 143810 61400 143866
rect 32606 143556 32998 143612
rect 33054 143556 33936 143612
rect 58240 143556 75348 143612
rect 75404 143556 75444 143612
rect 32658 143332 32802 143388
rect 32858 143332 33936 143388
rect 58240 143332 76020 143388
rect 76076 143332 76116 143388
rect 32658 143108 33054 143164
rect 33110 143108 33936 143164
rect 58240 143108 76692 143164
rect 76748 143108 76788 143164
rect 32658 142884 33306 142940
rect 33362 142884 33936 142940
rect 58240 142884 77364 142940
rect 77420 142884 77460 142940
rect 32658 142660 33558 142716
rect 33614 142660 33936 142716
rect 58240 142660 67284 142716
rect 67340 142660 67380 142716
rect 32658 142436 33810 142492
rect 33866 142436 33936 142492
rect 58240 142436 67956 142492
rect 68012 142436 68052 142492
rect 81144 142380 81270 146412
rect 81648 142380 81774 146412
rect 147212 146372 147252 146428
rect 147308 146372 313586 146428
rect 313642 146372 313682 146428
rect 149452 146250 149492 146306
rect 149548 146250 313334 146306
rect 313390 146250 313430 146306
rect 151692 146128 151732 146184
rect 151788 146128 313082 146184
rect 313138 146128 313178 146184
rect 153932 146006 153972 146062
rect 154028 146006 312830 146062
rect 312886 146006 312926 146062
rect 156172 145884 156212 145940
rect 156268 145884 312578 145940
rect 312634 145884 312674 145940
rect 158412 145762 158452 145818
rect 158508 145762 312326 145818
rect 312382 145762 312422 145818
rect 160652 145640 160692 145696
rect 160748 145640 312074 145696
rect 312130 145640 312170 145696
rect 163340 145518 163380 145574
rect 163436 145518 311822 145574
rect 311878 145518 311918 145574
rect 165580 145396 165620 145452
rect 165676 145396 311570 145452
rect 311626 145396 311666 145452
rect 167820 145274 167860 145330
rect 167916 145274 311318 145330
rect 311374 145274 311414 145330
rect 170060 145152 170100 145208
rect 170156 145152 311066 145208
rect 311122 145152 311162 145208
rect 82432 144978 83216 145040
rect 172300 145030 172340 145086
rect 172396 145030 310814 145086
rect 310870 145030 310910 145086
rect 82432 144633 82494 144978
rect 83152 144633 83216 144978
rect 174540 144908 174580 144964
rect 174636 144908 310562 144964
rect 310618 144908 310658 144964
rect 176780 144786 176820 144842
rect 176876 144786 310310 144842
rect 310366 144786 310406 144842
rect 179020 144664 179060 144720
rect 179116 144664 310058 144720
rect 310114 144664 310154 144720
rect 82432 144592 83216 144633
rect 181708 144542 181748 144598
rect 181804 144542 309806 144598
rect 309862 144542 309902 144598
rect 183948 144420 183988 144476
rect 184044 144420 309554 144476
rect 309610 144420 309650 144476
rect 186188 144298 186228 144354
rect 186284 144298 309302 144354
rect 309358 144298 309398 144354
rect 188428 144176 188468 144232
rect 188524 144176 309050 144232
rect 309106 144176 309146 144232
rect 190668 144054 190708 144110
rect 190764 144054 308798 144110
rect 308854 144054 308894 144110
rect 192908 143932 192948 143988
rect 193004 143932 308546 143988
rect 308602 143932 308642 143988
rect 195148 143810 195188 143866
rect 195244 143810 308294 143866
rect 308350 143810 308390 143866
rect 197388 143688 197428 143744
rect 197484 143688 308042 143744
rect 308098 143688 308138 143744
rect 117420 143566 117460 143622
rect 117516 143566 307790 143622
rect 307846 143566 307886 143622
rect 117644 143444 117684 143500
rect 117740 143444 307538 143500
rect 307594 143444 307634 143500
rect 117868 143322 117908 143378
rect 117964 143322 307286 143378
rect 307342 143322 307382 143378
rect 118092 143200 118132 143256
rect 118188 143200 307034 143256
rect 307090 143200 307130 143256
rect 118316 143078 118356 143134
rect 118412 143078 306782 143134
rect 306838 143078 306878 143134
rect 118540 142956 118580 143012
rect 118636 142956 306530 143012
rect 306586 142956 306626 143012
rect 118764 142834 118804 142890
rect 118860 142834 306278 142890
rect 306334 142834 306374 142890
rect 118988 142712 119028 142768
rect 119084 142712 306026 142768
rect 306082 142712 306122 142768
rect 126940 142590 126980 142646
rect 127036 142590 305774 142646
rect 305830 142590 305870 142646
rect 129180 142468 129220 142524
rect 129276 142468 305522 142524
rect 305578 142468 305618 142524
rect 58240 142212 68628 142268
rect 68684 142212 68724 142268
rect 81144 142254 81774 142380
rect 131420 142346 131460 142402
rect 131516 142346 305270 142402
rect 305326 142346 305366 142402
rect 133660 142224 133700 142280
rect 133756 142224 305018 142280
rect 305074 142224 305114 142280
rect 135900 142102 135940 142158
rect 135996 142102 304766 142158
rect 304822 142102 304862 142158
rect 58240 141988 69300 142044
rect 69356 141988 69396 142044
rect 138140 141980 138180 142036
rect 138236 141980 304514 142036
rect 304570 141980 304610 142036
rect 140380 141858 140420 141914
rect 140476 141858 304262 141914
rect 304318 141858 304358 141914
rect 58240 141764 69972 141820
rect 70028 141764 70068 141820
rect 142620 141736 142660 141792
rect 142716 141736 304010 141792
rect 304066 141736 304106 141792
rect 145308 141614 145348 141670
rect 145404 141614 303758 141670
rect 303814 141614 303854 141670
rect 58240 141540 70644 141596
rect 70700 141540 70740 141596
rect 147548 141492 147588 141548
rect 147644 141492 303506 141548
rect 303562 141492 303602 141548
rect 58240 141316 71316 141372
rect 71372 141316 71412 141372
rect 149788 141370 149828 141426
rect 149884 141370 303254 141426
rect 303310 141370 303350 141426
rect 152028 141248 152068 141304
rect 152124 141248 303002 141304
rect 303058 141248 303098 141304
rect 58240 141092 71988 141148
rect 72044 141092 72084 141148
rect 154268 141126 154308 141182
rect 154364 141126 302750 141182
rect 302806 141126 302846 141182
rect 156508 141004 156548 141060
rect 156604 141004 302498 141060
rect 302554 141004 302594 141060
rect 58240 140868 72660 140924
rect 72716 140868 72756 140924
rect 158748 140882 158788 140938
rect 158844 140882 302246 140938
rect 302302 140882 302342 140938
rect 160988 140760 161028 140816
rect 161084 140760 301994 140816
rect 302050 140760 302090 140816
rect 58240 140644 73332 140700
rect 73388 140644 73428 140700
rect 163676 140638 163716 140694
rect 163772 140638 301742 140694
rect 301798 140638 301838 140694
rect 165916 140516 165956 140572
rect 166012 140516 301490 140572
rect 301546 140516 301586 140572
rect 58240 140420 74004 140476
rect 74060 140420 74100 140476
rect 168156 140394 168196 140450
rect 168252 140394 301238 140450
rect 301294 140394 301334 140450
rect 170396 140272 170436 140328
rect 170492 140272 300986 140328
rect 301042 140272 301082 140328
rect 58240 140196 74676 140252
rect 74732 140196 74772 140252
rect 172636 140150 172676 140206
rect 172732 140150 300734 140206
rect 300790 140150 300830 140206
rect 174876 140028 174916 140084
rect 174972 140028 300482 140084
rect 300538 140028 300578 140084
rect 58240 139972 58548 140028
rect 58604 139972 59836 140028
rect 177116 139906 177156 139962
rect 177212 139906 300230 139962
rect 300286 139906 300326 139962
rect 58240 139748 78036 139804
rect 78092 139748 78132 139804
rect 179356 139784 179396 139840
rect 179452 139784 299978 139840
rect 300034 139784 300074 139840
rect 182044 139662 182084 139718
rect 182140 139662 299726 139718
rect 299782 139662 299822 139718
rect 58240 139524 78708 139580
rect 78764 139524 78804 139580
rect 184284 139540 184324 139596
rect 184380 139540 299474 139596
rect 299530 139540 299570 139596
rect 58240 139300 79380 139356
rect 79436 139300 79476 139356
rect 89152 139328 90832 139440
rect 186524 139418 186564 139474
rect 186620 139418 299222 139474
rect 299278 139418 299318 139474
rect 58240 139076 61908 139132
rect 61964 139076 62004 139132
rect 58240 138852 62580 138908
rect 62636 138852 62676 138908
rect 58240 138628 63252 138684
rect 63308 138628 63348 138684
rect 58240 138404 63924 138460
rect 63980 138404 64020 138460
rect 89152 138432 89264 139328
rect 90720 138432 90832 139328
rect 188764 139296 188804 139352
rect 188860 139296 298970 139352
rect 299026 139296 299066 139352
rect 191004 139174 191044 139230
rect 191100 139174 298718 139230
rect 298774 139174 298814 139230
rect 193244 139052 193284 139108
rect 193340 139052 298466 139108
rect 298522 139052 298562 139108
rect 195484 138930 195524 138986
rect 195580 138930 298214 138986
rect 298270 138930 298310 138986
rect 197724 138808 197764 138864
rect 197820 138808 297962 138864
rect 298018 138808 298058 138864
rect 125484 138686 125524 138742
rect 125580 138686 297710 138742
rect 297766 138686 297806 138742
rect 123580 138564 123620 138620
rect 123676 138564 297458 138620
rect 297514 138564 297554 138620
rect 125820 138442 125860 138498
rect 125916 138442 297206 138498
rect 297262 138442 297302 138498
rect 89152 138320 90832 138432
rect 117196 138320 117236 138376
rect 117292 138320 296954 138376
rect 297010 138320 297050 138376
rect 58240 138180 64596 138236
rect 64652 138180 64692 138236
rect 115852 138198 115892 138254
rect 115948 138198 296702 138254
rect 296758 138198 296798 138254
rect 116076 138076 116116 138132
rect 116172 138076 296450 138132
rect 296506 138076 296546 138132
rect 58240 137956 65268 138012
rect 65324 137956 65364 138012
rect 116524 137954 116564 138010
rect 116620 137954 296198 138010
rect 296254 137954 296294 138010
rect 116300 137832 116340 137888
rect 116396 137832 295946 137888
rect 296002 137832 296042 137888
rect 58240 137732 65940 137788
rect 65996 137732 66036 137788
rect 86958 137710 86968 137766
rect 87024 137710 295694 137766
rect 295750 137710 295771 137766
rect 58240 137508 66612 137564
rect 66668 137508 66708 137564
rect 58240 137284 58324 137340
rect 58380 137284 72548 137340
rect 72604 137284 72644 137340
rect 83626 137312 83636 137368
rect 83692 137312 124628 137368
rect 124684 137312 206990 137368
rect 207046 137312 207056 137368
rect 58240 137060 73220 137116
rect 73276 137060 73316 137116
rect 58240 136276 70532 136332
rect 70588 136276 70628 136332
rect 58240 136052 71204 136108
rect 71260 136052 71300 136108
rect 60858 135828 61488 135954
rect 60858 133560 60984 135828
rect 61362 133560 61488 135828
rect 60858 133434 61488 133560
rect 275800 133700 276600 133800
rect 275800 133100 275900 133700
rect 276500 133100 276600 133700
rect 275800 133000 276600 133100
rect 72188 132804 73196 132930
rect 72188 132174 72314 132804
rect 73070 132174 73196 132804
rect 72188 132048 73196 132174
rect 275800 132300 276600 132400
rect 66602 131908 66612 131964
rect 66668 131908 67172 131964
rect 67228 131908 67732 131964
rect 67788 131908 68852 131964
rect 68908 131908 69412 131964
rect 69468 131908 69972 131964
rect 70028 131908 70532 131964
rect 70588 131908 70598 131964
rect 275800 131700 275900 132300
rect 276500 131700 276600 132300
rect 58240 131572 71876 131628
rect 71932 131572 71972 131628
rect 275800 131600 276600 131700
rect 62622 131292 65772 131418
rect 62622 131040 62748 131292
rect 65646 131040 65772 131292
rect 62622 130914 65772 131040
rect 68941 130577 68964 130633
rect 69020 130577 86282 130633
rect 86338 130577 86363 130633
rect 59850 130511 60102 130536
rect 59850 130057 59875 130511
rect 60078 130057 60102 130511
rect 59850 130032 60102 130057
rect 61611 130477 61897 130534
rect 61611 130051 61634 130477
rect 61874 130051 61897 130477
rect 61611 130030 61897 130051
rect 62622 130410 65772 130536
rect 62622 130158 62748 130410
rect 65646 130158 65772 130410
rect 62622 130032 65772 130158
rect 58240 129780 69860 129836
rect 69916 129780 69956 129836
rect 202328 129379 202384 129410
rect 58240 128884 68964 128940
rect 69020 128884 69060 128940
rect 58240 128212 69188 128268
rect 69244 128212 69284 128268
rect 58240 127988 60340 128044
rect 60396 127988 60480 128044
rect 59724 127638 60228 127764
rect 59724 127386 59850 127638
rect 60102 127386 60228 127638
rect 59724 127260 60228 127386
rect 60984 127008 61992 127134
rect 60984 126630 61110 127008
rect 61866 126630 61992 127008
rect 60984 126504 61992 126630
rect 58240 126196 67396 126252
rect 67452 126196 67492 126252
rect 66528 124852 66612 124908
rect 66668 124852 81788 124908
rect 59024 124628 59114 124684
rect 59194 124628 81564 124684
rect 56268 124404 56308 124460
rect 56364 124404 73892 124460
rect 73948 124404 73988 124460
rect 53244 124180 53284 124236
rect 53340 124180 74564 124236
rect 74620 124180 74660 124236
rect 52684 123956 52724 124012
rect 52780 123956 75236 124012
rect 75292 123956 75332 124012
rect 52460 123732 52500 123788
rect 52556 123732 75908 123788
rect 75964 123732 76004 123788
rect 52236 123508 52276 123564
rect 52332 123508 77252 123564
rect 77308 123508 77348 123564
rect 52012 123284 52052 123340
rect 52108 123284 77924 123340
rect 77980 123284 78020 123340
rect 81508 123228 81564 124628
rect 81732 123452 81788 124852
rect 81732 123396 115220 123452
rect 115276 123396 115286 123452
rect 81508 123217 115388 123228
rect 81492 123161 115387 123217
rect 115443 123161 115467 123217
rect 51788 123060 51828 123116
rect 51884 123060 78596 123116
rect 78652 123060 78692 123116
rect 48876 122836 48916 122892
rect 48972 122836 79268 122892
rect 79324 122836 79364 122892
rect 44284 122612 44324 122668
rect 44380 122612 76580 122668
rect 76636 122612 76676 122668
rect 79676 122612 79716 122668
rect 79772 122612 113784 122668
rect 32504 122368 32550 122424
rect 32606 122368 66612 122424
rect 66668 122368 66708 122424
rect 79004 122388 79044 122444
rect 79100 122388 113560 122444
rect 78332 122164 78372 122220
rect 78428 122164 113336 122220
rect 77660 121940 77700 121996
rect 77756 121940 113112 121996
rect 70536 121716 70550 121772
rect 70606 121716 80500 121772
rect 80556 121716 80566 121772
rect 39320 121492 39360 121548
rect 39428 121492 74340 121548
rect 74396 121492 74436 121548
rect 39192 121268 39232 121324
rect 39300 121268 75012 121324
rect 75068 121268 75108 121324
rect 39064 121044 39104 121100
rect 39172 121044 75684 121100
rect 75740 121044 75780 121100
rect 38936 120820 38976 120876
rect 39044 120820 76356 120876
rect 76412 120820 76452 120876
rect 32550 119202 32606 119324
rect 32550 75674 32606 118958
rect 32550 75334 32606 75374
rect 32802 119202 32858 119324
rect 32802 75674 32858 118958
rect 32802 75334 32858 75374
rect 33054 119202 33110 119324
rect 33054 75674 33110 118958
rect 33054 75334 33110 75374
rect 33306 119202 33362 119324
rect 33306 75674 33362 118958
rect 33306 75334 33362 75374
rect 33558 119202 33614 119324
rect 33558 75674 33614 118958
rect 33558 75334 33614 75374
rect 33810 119202 33866 119324
rect 33810 75674 33866 118958
rect 113056 117996 113112 121940
rect 113280 118220 113336 122164
rect 113504 118444 113560 122388
rect 113728 118668 113784 122612
rect 113728 118612 118132 118668
rect 118188 118612 118228 118668
rect 113504 118388 117908 118444
rect 117964 118388 118004 118444
rect 113280 118164 117684 118220
rect 117740 118164 117780 118220
rect 113056 117940 117460 117996
rect 117516 117940 117556 117996
rect 34524 116046 35532 116172
rect 34524 114912 34650 116046
rect 35406 114912 35532 116046
rect 34524 114786 35532 114912
rect 90342 110880 90972 111006
rect 73458 110609 73710 110628
rect 73458 110390 73470 110609
rect 73693 110390 73710 110609
rect 58962 110054 59000 110110
rect 59056 110054 70980 110110
rect 71036 110054 71086 110110
rect 34309 109620 38682 109746
rect 34309 109085 37674 109620
rect 34309 101246 34333 109085
rect 34506 108612 37674 109085
rect 38556 108612 38682 109620
rect 73458 109620 73710 110390
rect 90342 110502 90468 110880
rect 90846 110502 90972 110880
rect 90342 110376 90972 110502
rect 103950 110376 107856 110502
rect 91350 109620 91854 109746
rect 73458 109368 86412 109620
rect 86640 109368 86656 109620
rect 66780 109116 67662 109242
rect 66780 108738 66906 109116
rect 67536 108738 67662 109116
rect 66780 108612 67662 108738
rect 91350 108738 91476 109620
rect 91728 108738 91854 109620
rect 91350 108612 91854 108738
rect 34506 108486 38682 108612
rect 70980 108500 71008 108556
rect 71450 108500 80836 108556
rect 80892 108500 80918 108556
rect 34506 101246 37303 108486
rect 37851 107984 37870 108040
rect 38167 107984 58324 108040
rect 58380 107984 58408 108040
rect 74214 107856 75222 107982
rect 37849 107648 37870 107704
rect 38167 107648 61486 107704
rect 61546 107648 61567 107704
rect 65772 107604 66654 107730
rect 59472 107352 60732 107478
rect 59472 106974 59598 107352
rect 60606 106974 60732 107352
rect 65772 107226 65898 107604
rect 66528 107226 66654 107604
rect 74214 107352 74340 107856
rect 75096 107352 75222 107856
rect 74214 107226 75222 107352
rect 92358 107856 93114 107982
rect 92358 107352 92484 107856
rect 92988 107352 93114 107856
rect 92358 107226 93114 107352
rect 65772 107100 66654 107226
rect 59472 106848 60732 106974
rect 77324 107084 103156 107140
rect 77324 106746 77380 107084
rect 77848 106755 77864 106907
rect 77932 106755 102081 106907
rect 102141 106755 102481 106907
rect 102541 106755 102551 106907
rect 73456 106690 73472 106746
rect 73528 106690 77380 106746
rect 39543 106453 39560 106605
rect 39628 106453 102281 106605
rect 102341 106453 102681 106605
rect 102741 106453 102760 106605
rect 103100 106508 103156 107084
rect 103100 106422 103156 106452
rect 103950 107100 104076 110376
rect 107730 107100 107856 110376
rect 103950 106852 107856 107100
rect 41172 106254 41220 106310
rect 41288 106254 59000 106310
rect 59056 106254 59094 106310
rect 62360 106198 62384 106254
rect 62658 106198 68450 106254
rect 68678 106198 68692 106254
rect 71628 106248 71652 106304
rect 71708 106248 77696 106304
rect 77764 106248 77777 106304
rect 103950 105588 105739 106852
rect 106057 105588 107856 106852
rect 34309 76576 37303 101246
rect 98784 84879 100010 85005
rect 100258 84934 101343 85005
rect 98784 82782 98910 84879
rect 99920 82782 100010 84879
rect 98784 82656 100010 82782
rect 100254 84884 101343 84934
rect 101591 84932 102630 85005
rect 100254 84879 101346 84884
rect 100254 82782 100344 84879
rect 101224 82782 101346 84879
rect 100254 82760 101346 82782
rect 100258 82710 101346 82760
rect 101590 84879 102630 84932
rect 102878 84914 104328 85005
rect 101590 82782 101680 84879
rect 102540 82782 102630 84879
rect 101590 82758 102630 82782
rect 100258 82656 101343 82710
rect 101591 82656 102630 82758
rect 102877 84879 104328 84914
rect 102877 82782 102967 84879
rect 104202 82782 104328 84879
rect 102877 82740 104328 82782
rect 102878 82656 104328 82740
rect 116300 81876 116340 81932
rect 116396 81876 119979 81932
rect 116524 80644 116564 80700
rect 116620 80644 119979 80700
rect 202328 78411 202384 129086
rect 202328 78097 202384 78126
rect 203084 129380 203140 129410
rect 203084 78404 203140 129075
rect 203084 78097 203140 78128
rect 203336 129385 203392 129410
rect 203336 78404 203392 129062
rect 203336 78097 203392 78128
rect 203588 129372 203644 129410
rect 203588 78404 203644 129064
rect 203588 78097 203644 78128
rect 203840 129370 203896 129410
rect 203840 78404 203896 129061
rect 203840 78097 203896 78128
rect 206990 120204 207046 120232
rect 206990 78624 207046 119700
rect 477200 79400 477800 79500
rect 477200 79000 477300 79400
rect 477700 79000 477800 79400
rect 477200 78900 477800 79000
rect 206990 78092 207046 78120
rect 477200 78400 477800 78500
rect 115643 77956 115668 78012
rect 115724 77956 119979 78012
rect 477200 78000 477300 78400
rect 477700 78000 477800 78400
rect 477200 77900 477800 78000
rect 201666 77344 207874 77417
rect 201639 77140 207898 77213
rect 201639 76936 207898 77009
rect 201639 76732 207898 76805
rect 201639 76528 207898 76601
rect 201639 76324 207898 76397
rect 472400 75600 478000 75800
rect 207589 75404 207645 75414
rect 33810 75334 33866 75374
rect 115658 75348 115668 75404
rect 115724 75348 122388 75404
rect 122444 75348 124404 75404
rect 124460 75348 128436 75404
rect 128492 75348 207589 75404
rect 207589 75338 207645 75348
rect 115839 74693 115849 74749
rect 115905 74693 126420 74749
rect 126476 74693 126486 74749
rect 135946 72828 140986 72954
rect 114597 72198 115227 72261
rect 113148 72072 114030 72198
rect 36236 71588 36288 71868
rect 36848 71588 112494 71868
rect 112570 71588 112598 71868
rect 113148 71442 113274 72072
rect 113904 71442 114030 72072
rect 113148 71316 114030 71442
rect 114597 71694 114660 72198
rect 115164 71694 115227 72198
rect 114597 71064 115227 71694
rect 135946 71442 136072 72828
rect 140860 71442 140986 72828
rect 135946 71316 140986 71442
rect 96894 70938 115227 71064
rect 96894 69426 97020 70938
rect 106218 70434 115227 70938
rect 106218 69426 106344 70434
rect 96894 69300 106344 69426
rect 208656 61768 208801 62370
rect 208656 61668 208801 61712
rect 213764 59885 213886 62364
rect 268380 61362 283248 61488
rect 268380 59472 268506 61362
rect 283122 59472 283248 61362
rect 472400 61200 472600 75600
rect 477800 61200 478000 75600
rect 472400 61000 478000 61200
rect 268380 59346 283248 59472
rect 213764 58937 213886 58998
rect 285200 58600 300000 58800
rect 34400 57600 36400 57800
rect 34400 43200 34600 57600
rect 36200 43200 36400 57600
rect 199000 53800 204646 54000
rect 199000 51600 199200 53800
rect 204464 51600 204646 53800
rect 199000 51400 204646 51600
rect 205266 53800 211000 54000
rect 205266 51600 205440 53800
rect 210800 51600 211000 53800
rect 285200 53400 285400 58600
rect 299800 53400 300000 58600
rect 285200 53200 300000 53400
rect 317800 52300 318600 52400
rect 317800 51700 317900 52300
rect 318500 51700 318600 52300
rect 317800 51600 318600 51700
rect 205266 51400 211000 51600
rect 317800 51100 318600 51200
rect 96138 50526 97603 50652
rect 96138 47754 96264 50526
rect 97476 47754 97603 50526
rect 96138 47628 97603 47754
rect 97872 50526 99412 50652
rect 97872 47754 97964 50526
rect 99320 47754 99412 50526
rect 97872 47628 99412 47754
rect 99669 50643 100639 50652
rect 101119 50646 101937 50652
rect 99669 50526 100640 50643
rect 99669 47754 99742 50526
rect 100567 47754 100640 50526
rect 99669 47660 100640 47754
rect 100893 50526 101937 50646
rect 102194 50627 103107 50652
rect 103364 50631 104748 50652
rect 102191 50526 103107 50627
rect 100893 47754 100966 50526
rect 101841 47754 101934 50526
rect 102191 47754 102284 50526
rect 103006 47754 103107 50526
rect 100893 47699 101937 47754
rect 99669 47628 100639 47660
rect 100896 47628 101937 47699
rect 102191 47695 103107 47754
rect 102194 47628 103107 47695
rect 103360 50526 104748 50631
rect 105005 50627 105917 50652
rect 103360 47754 103453 50526
rect 104649 47754 104748 50526
rect 103360 47628 104748 47754
rect 105003 50526 105917 50627
rect 105003 47754 105096 50526
rect 105822 47754 105917 50526
rect 105003 47695 105917 47754
rect 105005 47628 105917 47695
rect 106174 50526 107604 50652
rect 106174 47754 106276 50526
rect 107478 47754 107604 50526
rect 317800 50500 317900 51100
rect 318500 50500 318600 51100
rect 317800 50400 318600 50500
rect 106174 47628 107604 47754
rect 480400 45100 481200 45200
rect 480400 44500 480500 45100
rect 481100 44500 481200 45100
rect 480400 44400 481200 44500
rect 34400 43000 36400 43200
rect 480400 43700 481200 43800
rect 480400 43100 480500 43700
rect 481100 43100 481200 43700
rect 480400 43000 481200 43100
rect 231600 42200 246400 42400
rect 59700 41700 60500 41800
rect 59700 41100 59800 41700
rect 60400 41100 60500 41700
rect 59700 41000 60500 41100
rect 59700 40500 60500 40600
rect 59700 39900 59800 40500
rect 60400 39900 60500 40500
rect 59700 39800 60500 39900
rect 231600 37200 231800 42200
rect 246200 37200 246400 42200
rect 231600 37000 246400 37200
rect 102200 35400 117000 35600
rect 102200 33800 102400 35400
rect 116800 33800 117000 35400
rect 102200 33600 117000 33800
rect 300244 34969 300300 34979
rect 300244 33404 300300 34913
rect 300244 33338 300300 33348
<< via3 >>
rect 33600 366000 34600 380400
rect 332154 380250 332744 380778
rect 427400 374200 441800 375800
rect 444200 374200 458600 375800
rect 467000 374200 481400 375800
rect 470300 373000 470800 373500
rect 471500 373000 472000 373500
rect 63504 366912 64764 367542
rect 33600 349200 34600 363600
rect 320796 364604 322686 365486
rect 328600 364800 329200 365400
rect 328600 363400 329200 364000
rect 65394 360360 65646 360864
rect 66150 360360 66780 361620
rect 316890 360612 317646 360990
rect 63126 358092 63378 358470
rect 41076 356958 44604 357210
rect 60102 357084 62748 357336
rect 37800 337428 40068 338184
rect 49518 337428 51786 338184
rect 61992 337554 64260 338310
rect 322056 361872 323316 362502
rect 334600 360800 346000 362200
rect 326340 359226 329364 359982
rect 472600 349200 477800 363600
rect 410256 340578 411894 341712
rect 328230 340074 338814 340452
rect 33120 335888 33462 336226
rect 37800 334404 40068 335160
rect 49518 334530 51786 335286
rect 61992 334404 64260 335160
rect 37674 315378 38682 315630
rect 52668 315504 54054 315756
rect 63756 315378 65016 315630
rect 35154 312984 35910 313488
rect 38413 313329 38578 313604
rect 41744 313357 41962 313623
rect 42840 312858 43218 313614
rect 44030 313428 44407 313687
rect 45467 313339 45631 313601
rect 48779 313364 49011 313634
rect 60354 313110 61236 313362
rect 64512 312480 65394 312732
rect 50283 312160 50882 312393
rect 60354 311472 61236 311724
rect 68670 310968 69426 311220
rect 42840 310338 43218 310842
rect 50022 310338 50400 310842
rect 64386 310716 65520 310842
rect 57903 310206 58105 310424
rect 50652 309078 51282 309582
rect 58590 308952 58842 309582
rect 32550 308528 32810 308767
rect 38386 308528 38625 308767
rect 45418 308528 45657 308767
rect 33150 308123 33410 308296
rect 59346 307062 61362 307692
rect 57960 287910 60354 288162
rect 49186 283673 50234 283951
rect 54858 283680 55884 283944
rect 34950 281649 35210 282082
rect 33739 254062 33994 257206
rect 35550 248888 35810 249475
rect 58590 247086 59220 247968
rect 60228 245448 60858 246330
rect 63882 243936 64638 244692
rect 67284 242298 67914 243180
rect 65764 241290 66898 241794
rect 34339 237262 34594 240406
rect 49770 239778 51660 239904
rect 64857 238630 65097 239346
rect 34950 237449 35210 237882
rect 66402 232596 66654 233604
rect 72450 228690 73584 229320
rect 65394 225792 66528 226674
rect 33176 219357 33382 223223
rect 72954 208656 73584 209538
rect 79331 206980 79685 207942
rect 34939 203662 35194 206806
rect 35550 205288 35810 205875
rect 74345 205038 74614 205722
rect 73206 199710 73710 200970
rect 33750 198886 34010 199085
rect 32550 198151 32810 198350
rect 36150 197377 36410 197670
rect 49829 196869 51830 197117
rect 34950 194649 35210 195082
rect 35539 186862 35794 190006
rect 66150 189252 66780 190008
rect 70812 198094 71316 198850
rect 69048 192402 69552 193032
rect 65772 183078 66906 184212
rect 36139 170062 36394 173206
rect 73332 166446 74088 167202
rect 79506 164178 79884 165312
rect 35550 162488 35810 163075
rect 80892 161532 81522 162036
rect 70964 156500 71720 156752
rect 36739 153262 36994 156406
rect 72072 156492 72828 156744
rect 51408 152838 52794 153468
rect 321100 149336 321500 149736
rect 321100 148336 321500 148736
rect 81270 142380 81648 146412
rect 82494 144633 83152 144978
rect 89264 138432 90720 139328
rect 60984 133560 61362 135828
rect 275900 133100 276500 133700
rect 72314 132174 73070 132804
rect 275900 131700 276500 132300
rect 62748 131040 65646 131292
rect 59875 130057 60078 130511
rect 61634 130051 61874 130477
rect 62748 130158 65646 130410
rect 59850 127386 60102 127638
rect 61110 126630 61866 127008
rect 34650 114912 35406 116046
rect 73470 110390 73693 110609
rect 37674 108612 38556 109620
rect 90468 110502 90846 110880
rect 66906 108738 67536 109116
rect 91476 108738 91728 109620
rect 59598 106974 60606 107352
rect 65898 107226 66528 107604
rect 74340 107352 75096 107856
rect 92484 107352 92988 107856
rect 104076 107100 107730 110376
rect 98910 82782 99920 84879
rect 100344 82782 101224 84879
rect 101680 82782 102540 84879
rect 102967 82782 104202 84879
rect 477300 79000 477700 79400
rect 477300 78000 477700 78400
rect 36288 71588 36848 71868
rect 113274 71442 113904 72072
rect 136072 71442 140860 72828
rect 97020 69426 106218 70938
rect 268506 59472 283122 61362
rect 472600 61200 477800 75600
rect 34600 43200 36200 57600
rect 199200 51600 204464 53800
rect 205440 51600 210800 53800
rect 285400 53400 299800 58600
rect 317900 51700 318500 52300
rect 96264 47754 97476 50526
rect 97964 47754 99320 50526
rect 99742 47754 100567 50526
rect 100966 47754 101841 50526
rect 102284 47754 103006 50526
rect 103453 47754 104649 50526
rect 105096 47754 105822 50526
rect 106276 47754 107478 50526
rect 317900 50500 318500 51100
rect 480500 44500 481100 45100
rect 480500 43100 481100 43700
rect 59800 41100 60400 41700
rect 59800 39900 60400 40500
rect 231800 37200 246200 42200
rect 102400 33800 116800 35400
<< metal4 >>
rect 332100 380778 332806 380830
rect 33400 380400 34800 380600
rect 33400 366000 33600 380400
rect 34600 366000 34800 380400
rect 332100 380250 332154 380778
rect 332744 380250 332806 380778
rect 332100 380188 332806 380250
rect 427200 375984 442000 376000
rect 413784 375800 442000 375984
rect 413784 374724 427400 375800
rect 413770 374200 427400 374724
rect 441800 374200 442000 375800
rect 413770 374000 442000 374200
rect 444000 375800 458800 376000
rect 444000 374200 444200 375800
rect 458600 374200 458800 375800
rect 444000 374000 447000 374200
rect 452600 374000 458800 374200
rect 466800 375800 481600 376000
rect 466800 374200 467000 375800
rect 481400 374200 481600 375800
rect 466800 374000 481600 374200
rect 33400 365800 34800 366000
rect 40950 368424 44730 368550
rect 40950 366786 41076 368424
rect 44604 366786 44730 368424
rect 33400 363600 34800 363800
rect 33400 349200 33600 363600
rect 34600 349200 34800 363600
rect 40950 357210 44730 366786
rect 40950 356958 41076 357210
rect 44604 356958 44730 357210
rect 59976 368046 62874 368172
rect 59976 366786 60102 368046
rect 62748 366786 62874 368046
rect 63378 367542 64890 367668
rect 63378 366912 63504 367542
rect 64764 366912 64890 367542
rect 63378 366786 64890 366912
rect 59976 357336 62874 366786
rect 320670 365486 322812 365612
rect 320670 364604 320796 365486
rect 322686 364604 322812 365486
rect 328500 365400 329300 365500
rect 328500 364800 328600 365400
rect 329200 364800 329300 365400
rect 328500 364700 329300 364800
rect 320670 364478 322812 364604
rect 328500 364000 329300 364100
rect 328500 363400 328600 364000
rect 329200 363400 329300 364000
rect 328500 363300 329300 363400
rect 326214 362880 329490 363006
rect 321930 362502 323442 362628
rect 321930 361872 322056 362502
rect 323316 361872 323442 362502
rect 321930 361746 323442 361872
rect 66024 361620 66906 361746
rect 65268 360864 65772 360990
rect 65268 360360 65394 360864
rect 65646 360360 65772 360864
rect 63000 358470 63504 358596
rect 63000 358092 63126 358470
rect 63378 358092 63504 358470
rect 63000 357966 63504 358092
rect 65268 358470 65772 360360
rect 66024 360360 66150 361620
rect 66780 360360 66906 361620
rect 326214 361242 326340 362880
rect 329364 361242 329490 362880
rect 66024 360234 66906 360360
rect 316764 360990 317898 361116
rect 316764 360612 316890 360990
rect 317646 360612 317898 360990
rect 65268 357714 65394 358470
rect 65646 357714 65772 358470
rect 65268 357588 65772 357714
rect 59976 357084 60102 357336
rect 62748 357084 62874 357336
rect 59976 356958 62874 357084
rect 40950 356832 44730 356958
rect 33400 349000 34800 349200
rect 316764 341712 317898 360612
rect 326214 359982 329490 361242
rect 334400 362200 346200 362400
rect 334400 360800 334600 362200
rect 346000 360800 346200 362200
rect 334400 360600 346200 360800
rect 326214 359226 326340 359982
rect 329364 359226 329490 359982
rect 326214 359100 329490 359226
rect 413770 341838 416416 374000
rect 470200 373500 470900 373600
rect 470200 373000 470300 373500
rect 470800 373000 470900 373500
rect 470200 372900 470900 373000
rect 471400 373500 472100 373600
rect 471400 373000 471500 373500
rect 472000 373000 472100 373500
rect 471400 372900 472100 373000
rect 472400 363600 478000 363800
rect 472400 349200 472600 363600
rect 477800 349200 478000 363600
rect 472400 349000 478000 349200
rect 410130 341712 416416 341838
rect 316764 340578 410256 341712
rect 411894 340578 416416 341712
rect 316764 340452 416416 340578
rect 316764 340074 328230 340452
rect 338814 340074 416367 340452
rect 316764 339696 416367 340074
rect 61866 338310 64386 338436
rect 37674 338184 40194 338310
rect 37674 337428 37800 338184
rect 40068 337428 40194 338184
rect 37674 336798 40194 337428
rect 33078 336226 33506 336260
rect 33078 335888 33120 336226
rect 33462 336144 33506 336226
rect 37674 336144 37800 336798
rect 33462 335980 37800 336144
rect 33462 335888 33506 335980
rect 33078 335846 33506 335888
rect 37674 335916 37800 335980
rect 40068 335916 40194 336798
rect 37674 335160 40194 335916
rect 37674 334404 37800 335160
rect 40068 334404 40194 335160
rect 49392 338184 51912 338310
rect 49392 337428 49518 338184
rect 51786 337428 51912 338184
rect 49392 336798 51912 337428
rect 49392 335916 49518 336798
rect 51786 335916 51912 336798
rect 49392 335286 51912 335916
rect 49392 334530 49518 335286
rect 51786 334530 51912 335286
rect 49392 334404 51912 334530
rect 61866 337554 61992 338310
rect 64260 337554 64386 338310
rect 61866 336798 64386 337554
rect 61866 335916 61992 336798
rect 64260 335916 64386 336798
rect 61866 335160 64386 335916
rect 61866 334404 61992 335160
rect 64260 334404 64386 335160
rect 37674 334278 40194 334404
rect 61866 334278 64386 334404
rect 328130 328600 329030 338794
rect 328130 323200 328200 328600
rect 329000 323200 329030 328600
rect 328130 316468 329030 323200
rect 329158 336200 330006 338794
rect 329158 330800 329300 336200
rect 329900 330800 330006 336200
rect 329158 316468 330006 330800
rect 330126 328600 330386 338794
rect 330126 323200 330200 328600
rect 330300 323200 330386 328600
rect 330126 316468 330386 323200
rect 330506 336200 330766 338794
rect 330506 330800 330600 336200
rect 330700 330800 330766 336200
rect 330506 316468 330766 330800
rect 330886 336200 331408 338794
rect 330886 330800 331000 336200
rect 331300 330800 331408 336200
rect 330886 316468 331408 330800
rect 331528 328600 332676 338794
rect 331528 323200 331600 328600
rect 332600 323200 332676 328600
rect 331528 316468 332676 323200
rect 332796 336200 333526 338794
rect 332796 330800 332900 336200
rect 333400 330800 333526 336200
rect 332796 316468 333526 330800
rect 333646 328600 334150 338794
rect 333646 323200 333700 328600
rect 334000 323200 334150 328600
rect 333646 316468 334150 323200
rect 334270 336200 334530 338794
rect 334270 330800 334300 336200
rect 334400 330800 334530 336200
rect 334270 316468 334530 330800
rect 334650 336200 335172 338794
rect 334650 330800 334700 336200
rect 335000 330800 335172 336200
rect 334650 316468 335172 330800
rect 335292 328600 336440 338794
rect 335292 323200 335400 328600
rect 336400 323200 336440 328600
rect 335292 316468 336440 323200
rect 336560 336200 337290 338794
rect 336560 330800 336700 336200
rect 337200 330800 337290 336200
rect 336560 316468 337290 330800
rect 337410 328600 337914 338794
rect 337410 323200 337500 328600
rect 337800 323200 337914 328600
rect 337410 316468 337914 323200
rect 338034 336200 338294 338794
rect 338034 330800 338100 336200
rect 338200 330800 338294 336200
rect 338034 316468 338294 330800
rect 338414 336200 338936 338794
rect 338414 330800 338500 336200
rect 338800 330800 338936 336200
rect 338414 316468 338936 330800
rect 339056 328600 340204 338794
rect 339056 323200 339200 328600
rect 340200 323200 340204 328600
rect 339056 316468 340204 323200
rect 340324 336200 341054 338794
rect 340324 330800 340500 336200
rect 341000 330800 341054 336200
rect 340324 316468 341054 330800
rect 341174 328600 341678 338794
rect 341174 323200 341300 328600
rect 341600 323200 341678 328600
rect 341174 316468 341678 323200
rect 341798 336200 342058 338794
rect 341798 330800 341900 336200
rect 342000 330800 342058 336200
rect 341798 316468 342058 330800
rect 342178 336200 342700 338794
rect 342178 330800 342300 336200
rect 342600 330800 342700 336200
rect 342178 316468 342700 330800
rect 342820 328600 343968 338794
rect 342820 323200 342900 328600
rect 343900 323200 343968 328600
rect 342820 316468 343968 323200
rect 344088 336200 344818 338794
rect 344088 330800 344200 336200
rect 344700 330800 344818 336200
rect 344088 316468 344818 330800
rect 344938 328600 345442 338794
rect 344938 323200 345000 328600
rect 345300 323200 345442 328600
rect 344938 316468 345442 323200
rect 345562 336200 345822 338794
rect 345562 330800 345600 336200
rect 345700 330800 345822 336200
rect 345562 316468 345822 330800
rect 345942 336200 346464 338794
rect 345942 330800 346100 336200
rect 346400 330800 346464 336200
rect 345942 316468 346464 330800
rect 346584 328600 347732 338794
rect 346584 323200 346700 328600
rect 347700 323200 347732 328600
rect 346584 316468 347732 323200
rect 347852 336200 348582 338794
rect 347852 330800 348000 336200
rect 348500 330800 348582 336200
rect 347852 316468 348582 330800
rect 348702 328600 349206 338794
rect 348702 323200 348800 328600
rect 349100 323200 349206 328600
rect 348702 316468 349206 323200
rect 349326 336200 349586 338794
rect 349326 330800 349400 336200
rect 349500 330800 349586 336200
rect 349326 316468 349586 330800
rect 349706 336200 350228 338794
rect 349706 330800 349800 336200
rect 350100 330800 350228 336200
rect 349706 316468 350228 330800
rect 350348 328600 351496 338794
rect 350348 323200 350400 328600
rect 351400 323200 351496 328600
rect 350348 316468 351496 323200
rect 351616 336200 352346 338794
rect 351616 330800 351700 336200
rect 352200 330800 352346 336200
rect 351616 316468 352346 330800
rect 352466 328600 352970 338794
rect 352466 323200 352600 328600
rect 352900 323200 352970 328600
rect 352466 316468 352970 323200
rect 353090 336200 353350 338794
rect 353090 330800 353200 336200
rect 353300 330800 353350 336200
rect 353090 316468 353350 330800
rect 353470 336200 353992 338794
rect 353470 330800 353600 336200
rect 353900 330800 353992 336200
rect 353470 316468 353992 330800
rect 354112 328600 355260 338794
rect 354112 323200 354200 328600
rect 355200 323200 355260 328600
rect 354112 316468 355260 323200
rect 355380 336200 356110 338794
rect 355380 330800 355500 336200
rect 356000 330800 356110 336200
rect 355380 316468 356110 330800
rect 356230 328600 356734 338794
rect 356230 323200 356300 328600
rect 356600 323200 356734 328600
rect 356230 316468 356734 323200
rect 356854 336200 357114 338794
rect 356854 330800 356900 336200
rect 357000 330800 357114 336200
rect 356854 316468 357114 330800
rect 357234 336200 357756 338794
rect 357234 330800 357300 336200
rect 357600 330800 357756 336200
rect 357234 316468 357756 330800
rect 357876 328600 359024 338794
rect 357876 323200 358000 328600
rect 359000 323200 359024 328600
rect 357876 316468 359024 323200
rect 359144 336200 359874 338794
rect 359144 330800 359300 336200
rect 359800 330800 359874 336200
rect 359144 316468 359874 330800
rect 359994 328600 360498 338794
rect 359994 323200 360100 328600
rect 360400 323200 360498 328600
rect 359994 316468 360498 323200
rect 360618 336200 360878 338794
rect 360618 330800 360700 336200
rect 360800 330800 360878 336200
rect 360618 316468 360878 330800
rect 360998 336200 361520 338794
rect 360998 330800 361100 336200
rect 361400 330800 361520 336200
rect 360998 316468 361520 330800
rect 361640 328600 362788 338794
rect 361640 323200 361700 328600
rect 362700 323200 362788 328600
rect 361640 316468 362788 323200
rect 362908 336200 363638 338794
rect 362908 330800 363000 336200
rect 363500 330800 363638 336200
rect 362908 316468 363638 330800
rect 363758 328600 364262 338794
rect 363758 323200 363900 328600
rect 364200 323200 364262 328600
rect 363758 316468 364262 323200
rect 364382 336200 364642 338794
rect 364382 330800 364500 336200
rect 364600 330800 364642 336200
rect 364382 316468 364642 330800
rect 364762 336200 365284 338794
rect 364762 330800 364900 336200
rect 365200 330800 365284 336200
rect 364762 316468 365284 330800
rect 365404 328600 366552 338794
rect 365404 323200 365500 328600
rect 366500 323200 366552 328600
rect 365404 316468 366552 323200
rect 366672 336200 367402 338794
rect 366672 330800 366800 336200
rect 367300 330800 367402 336200
rect 366672 316468 367402 330800
rect 367522 328600 368026 338794
rect 367522 323200 367600 328600
rect 367900 323200 368026 328600
rect 367522 316468 368026 323200
rect 368146 336200 368406 338794
rect 368146 330800 368200 336200
rect 368300 330800 368406 336200
rect 368146 316468 368406 330800
rect 368526 336200 369048 338794
rect 368526 330800 368600 336200
rect 368900 330800 369048 336200
rect 368526 316468 369048 330800
rect 369168 328600 370316 338794
rect 369168 323200 369200 328600
rect 370200 323200 370316 328600
rect 369168 316468 370316 323200
rect 370436 336200 371166 338794
rect 370436 330800 370600 336200
rect 371100 330800 371166 336200
rect 370436 316468 371166 330800
rect 371286 328600 371790 338794
rect 371286 323200 371400 328600
rect 371700 323200 371790 328600
rect 371286 316468 371790 323200
rect 371910 336200 372170 338794
rect 371910 330800 372000 336200
rect 372100 330800 372170 336200
rect 371910 316468 372170 330800
rect 372290 336200 372812 338794
rect 372290 330800 372400 336200
rect 372700 330800 372812 336200
rect 372290 316468 372812 330800
rect 372932 328600 374080 338794
rect 372932 323200 373000 328600
rect 374000 323200 374080 328600
rect 372932 316468 374080 323200
rect 374200 336200 374930 338794
rect 374200 330800 374300 336200
rect 374800 330800 374930 336200
rect 374200 316468 374930 330800
rect 375050 328600 375554 338794
rect 375050 323200 375100 328600
rect 375400 323200 375554 328600
rect 375050 316468 375554 323200
rect 375674 336200 375934 338794
rect 375674 330800 375800 336200
rect 375900 330800 375934 336200
rect 375674 316468 375934 330800
rect 376054 336200 376576 338794
rect 376054 330800 376200 336200
rect 376500 330800 376576 336200
rect 376054 316468 376576 330800
rect 376696 328600 377844 338794
rect 376696 323200 376800 328600
rect 377800 323200 377844 328600
rect 376696 316468 377844 323200
rect 377964 336200 378694 338794
rect 377964 330800 378100 336200
rect 378600 330800 378694 336200
rect 377964 316468 378694 330800
rect 378814 328600 379318 338794
rect 378814 323200 378900 328600
rect 379200 323200 379318 328600
rect 378814 316468 379318 323200
rect 379438 336200 379698 338794
rect 379438 330800 379500 336200
rect 379600 330800 379698 336200
rect 379438 316468 379698 330800
rect 379818 336200 380340 338794
rect 379818 330800 379900 336200
rect 380200 330800 380340 336200
rect 379818 316468 380340 330800
rect 380460 328600 381608 338794
rect 380460 323200 380600 328600
rect 381600 323200 381608 328600
rect 380460 316468 381608 323200
rect 381728 336200 382458 338794
rect 381728 330800 381800 336200
rect 382300 330800 382458 336200
rect 381728 316468 382458 330800
rect 382578 328600 383082 338794
rect 382578 323200 382700 328600
rect 383000 323200 383082 328600
rect 382578 316468 383082 323200
rect 383202 336200 383462 338794
rect 383202 330800 383300 336200
rect 383400 330800 383462 336200
rect 383202 316468 383462 330800
rect 383582 336200 384104 338794
rect 383582 330800 383700 336200
rect 384000 330800 384104 336200
rect 383582 316468 384104 330800
rect 384224 328600 385372 338794
rect 384224 323200 384300 328600
rect 385300 323200 385372 328600
rect 384224 316468 385372 323200
rect 385492 336200 386222 338794
rect 385492 330800 385600 336200
rect 386100 330800 386222 336200
rect 385492 316468 386222 330800
rect 386342 328600 386846 338794
rect 386342 323200 386400 328600
rect 386700 323200 386846 328600
rect 386342 316468 386846 323200
rect 386966 336200 387226 338794
rect 386966 330800 387100 336200
rect 387200 330800 387226 336200
rect 386966 316468 387226 330800
rect 387346 336200 387868 338794
rect 387346 330800 387500 336200
rect 387800 330800 387868 336200
rect 387346 316468 387868 330800
rect 387988 328600 389136 338794
rect 387988 323200 388100 328600
rect 389100 323200 389136 328600
rect 387988 316468 389136 323200
rect 389256 336200 389986 338794
rect 389256 330800 389400 336200
rect 389900 330800 389986 336200
rect 389256 316468 389986 330800
rect 390106 328600 390610 338794
rect 390106 323200 390200 328600
rect 390500 323200 390610 328600
rect 390106 316468 390610 323200
rect 390730 336200 391070 338794
rect 390730 330800 390800 336200
rect 391000 330800 391070 336200
rect 390730 316468 391070 330800
rect 391191 328600 391843 338794
rect 391191 323200 391300 328600
rect 391700 323200 391843 328600
rect 391191 316468 391843 323200
rect 392135 336200 392641 338794
rect 392135 330800 392200 336200
rect 392500 330800 392641 336200
rect 392135 316468 392641 330800
rect 392761 328600 394057 338794
rect 392761 323200 392800 328600
rect 393800 323200 394057 328600
rect 392761 316468 394057 323200
rect 394260 336200 395910 338794
rect 394260 330800 394300 336200
rect 395800 330800 395910 336200
rect 394260 316468 395910 330800
rect 396034 328600 396480 338794
rect 396034 323200 396100 328600
rect 396400 323200 396480 328600
rect 396034 316468 396480 323200
rect 396668 336200 397866 338794
rect 396668 330800 396800 336200
rect 397800 330800 397866 336200
rect 396668 316468 397866 330800
rect 398068 328600 400054 338794
rect 398068 323200 398200 328600
rect 400000 323200 400054 328600
rect 398068 316468 400054 323200
rect 400465 336200 401953 338794
rect 400465 330800 400600 336200
rect 401800 330800 401953 336200
rect 400465 316468 401953 330800
rect 402200 328600 403368 338794
rect 402200 323200 402300 328600
rect 403300 323200 403368 328600
rect 402200 316468 403368 323200
rect 403507 328600 404631 338794
rect 403507 323200 403600 328600
rect 404600 323200 404631 328600
rect 403507 316468 404631 323200
rect 404761 336200 405445 338794
rect 404761 330800 404900 336200
rect 405400 330800 405445 336200
rect 404761 316468 405445 330800
rect 405585 328600 406309 338794
rect 405585 323200 405700 328600
rect 406200 323200 406309 328600
rect 405585 316468 406309 323200
rect 406429 336200 406689 338794
rect 406429 330800 406500 336200
rect 406600 330800 406689 336200
rect 406429 316468 406689 330800
rect 406809 336200 407331 338794
rect 406809 330800 406900 336200
rect 407300 330800 407331 336200
rect 406809 316468 407331 330800
rect 407451 328600 408599 338794
rect 407451 323200 407500 328600
rect 408500 323200 408599 328600
rect 407451 316468 408599 323200
rect 408719 336200 409449 338794
rect 408719 330800 408800 336200
rect 409300 330800 409449 336200
rect 408719 316468 409449 330800
rect 409569 328600 410073 338794
rect 409569 323200 409700 328600
rect 410000 323200 410073 328600
rect 409569 316468 410073 323200
rect 410193 336200 410453 338794
rect 410193 330800 410300 336200
rect 410400 330800 410453 336200
rect 410193 316468 410453 330800
rect 410573 336200 411095 338794
rect 410573 330800 410700 336200
rect 411000 330800 411095 336200
rect 410573 316468 411095 330800
rect 411215 328600 412363 338794
rect 411215 323200 411300 328600
rect 412300 323200 412363 328600
rect 411215 316468 412363 323200
rect 412483 336200 413213 338794
rect 412483 330800 412600 336200
rect 413100 330800 413213 336200
rect 412483 316468 413213 330800
rect 413333 328600 413837 338794
rect 413333 323200 413400 328600
rect 413700 323200 413837 328600
rect 413333 316468 413837 323200
rect 413957 336200 414217 338794
rect 413957 330800 414000 336200
rect 414100 330800 414217 336200
rect 413957 316468 414217 330800
rect 414337 336200 414859 338794
rect 414337 330800 414400 336200
rect 414700 330800 414859 336200
rect 414337 316468 414859 330800
rect 414979 328600 416127 338794
rect 414979 323200 415100 328600
rect 416100 323200 416127 328600
rect 414979 316468 416127 323200
rect 416247 336200 416977 338794
rect 416247 330800 416400 336200
rect 416900 330800 416977 336200
rect 416247 316468 416977 330800
rect 417097 328600 417601 338794
rect 417097 323200 417200 328600
rect 417500 323200 417601 328600
rect 417097 316468 417601 323200
rect 417721 336200 417981 338794
rect 417721 330800 417800 336200
rect 417900 330800 417981 336200
rect 417721 316468 417981 330800
rect 418101 336200 418623 338794
rect 418101 330800 418200 336200
rect 418500 330800 418623 336200
rect 418101 316468 418623 330800
rect 418743 328600 419891 338794
rect 418743 323200 418800 328600
rect 419800 323200 419891 328600
rect 418743 316468 419891 323200
rect 420011 336200 420741 338794
rect 420011 330800 420100 336200
rect 420600 330800 420741 336200
rect 420011 316468 420741 330800
rect 420861 328600 421365 338794
rect 420861 323200 420900 328600
rect 421200 323200 421365 328600
rect 420861 316468 421365 323200
rect 421485 336200 421745 338794
rect 421485 330800 421600 336200
rect 421700 330800 421745 336200
rect 421485 316468 421745 330800
rect 421865 336200 422387 338794
rect 421865 330800 422000 336200
rect 422300 330800 422387 336200
rect 421865 316468 422387 330800
rect 422507 328600 423655 338794
rect 422507 323200 422600 328600
rect 423600 323200 423655 328600
rect 422507 316468 423655 323200
rect 423775 336200 424505 338794
rect 423775 330800 423900 336200
rect 424400 330800 424505 336200
rect 423775 316468 424505 330800
rect 424625 328600 425129 338794
rect 424625 323200 424700 328600
rect 425000 323200 425129 328600
rect 424625 316468 425129 323200
rect 425249 336200 425509 338794
rect 425249 330800 425300 336200
rect 425400 330800 425509 336200
rect 425249 316468 425509 330800
rect 425629 336200 426151 338794
rect 425629 330800 425700 336200
rect 426000 330800 426151 336200
rect 425629 316468 426151 330800
rect 426271 328600 427419 338794
rect 426271 323200 426400 328600
rect 427400 323200 427419 328600
rect 426271 316468 427419 323200
rect 427539 336200 428269 338794
rect 427539 330800 427600 336200
rect 428100 330800 428269 336200
rect 427539 316468 428269 330800
rect 428389 328600 428893 338794
rect 428389 323200 428500 328600
rect 428800 323200 428893 328600
rect 428389 316468 428893 323200
rect 429013 336200 429273 338794
rect 429013 330800 429100 336200
rect 429200 330800 429273 336200
rect 429013 316468 429273 330800
rect 429393 336200 429915 338794
rect 429393 330800 429500 336200
rect 429800 330800 429915 336200
rect 429393 316468 429915 330800
rect 430035 328600 431183 338794
rect 430035 323200 430100 328600
rect 431100 323200 431183 328600
rect 430035 316468 431183 323200
rect 431303 336200 432033 338794
rect 431303 330800 431400 336200
rect 431900 330800 432033 336200
rect 431303 316468 432033 330800
rect 432153 328600 432657 338794
rect 432153 323200 432300 328600
rect 432600 323200 432657 328600
rect 432153 316468 432657 323200
rect 432777 336200 433037 338794
rect 432777 330800 432800 336200
rect 432900 330800 433037 336200
rect 432777 316468 433037 330800
rect 433157 336200 433679 338794
rect 433157 330800 433300 336200
rect 433600 330800 433679 336200
rect 433157 316468 433679 330800
rect 433799 328600 434947 338794
rect 433799 323200 433900 328600
rect 434900 323200 434947 328600
rect 433799 316468 434947 323200
rect 435067 336200 435797 338794
rect 435067 330800 435200 336200
rect 435700 330800 435797 336200
rect 435067 316468 435797 330800
rect 435917 328600 436421 338794
rect 435917 323200 436000 328600
rect 436300 323200 436421 328600
rect 435917 316468 436421 323200
rect 436541 336200 436801 338794
rect 436541 330800 436600 336200
rect 436700 330800 436801 336200
rect 436541 316468 436801 330800
rect 436921 336200 437443 338794
rect 436921 330800 437000 336200
rect 437300 330800 437443 336200
rect 436921 316468 437443 330800
rect 437563 328600 438711 338794
rect 437563 323200 437600 328600
rect 438600 323200 438711 328600
rect 437563 316468 438711 323200
rect 438831 336200 439561 338794
rect 438831 330800 438900 336200
rect 439400 330800 439561 336200
rect 438831 316468 439561 330800
rect 439681 328600 440185 338794
rect 439681 323200 439800 328600
rect 440100 323200 440185 328600
rect 439681 316468 440185 323200
rect 440305 336200 440565 338794
rect 440305 330800 440400 336200
rect 440500 330800 440565 336200
rect 440305 316468 440565 330800
rect 440685 336200 441207 338794
rect 440685 330800 440800 336200
rect 441100 330800 441207 336200
rect 440685 316468 441207 330800
rect 441327 328600 442475 338794
rect 441327 323200 441400 328600
rect 442400 323200 442475 328600
rect 441327 316468 442475 323200
rect 442595 336200 443325 338794
rect 442595 330800 442700 336200
rect 443200 330800 443325 336200
rect 442595 316468 443325 330800
rect 443445 328600 443949 338794
rect 443445 323200 443500 328600
rect 443800 323200 443949 328600
rect 443445 316468 443949 323200
rect 444069 336200 444329 338794
rect 444069 330800 444100 336200
rect 444200 330800 444329 336200
rect 444069 316468 444329 330800
rect 444449 336200 444971 338794
rect 444449 330800 444600 336200
rect 444900 330800 444971 336200
rect 444449 316468 444971 330800
rect 445091 328600 446239 338794
rect 445091 323200 445200 328600
rect 446200 323200 446239 328600
rect 445091 316468 446239 323200
rect 446359 336200 447089 338794
rect 446359 330800 446500 336200
rect 447000 330800 447089 336200
rect 446359 316468 447089 330800
rect 447209 328600 447713 338794
rect 447209 323200 447300 328600
rect 447600 323200 447713 328600
rect 447209 316468 447713 323200
rect 447833 336200 448093 338794
rect 447833 330800 447900 336200
rect 448000 330800 448093 336200
rect 447833 316468 448093 330800
rect 448213 336200 448735 338794
rect 448213 330800 448300 336200
rect 448600 330800 448735 336200
rect 448213 316468 448735 330800
rect 448855 328600 450003 338794
rect 448855 323200 448900 328600
rect 449900 323200 450003 328600
rect 448855 316468 450003 323200
rect 450123 336200 450853 338794
rect 450123 330800 450200 336200
rect 450700 330800 450853 336200
rect 450123 316468 450853 330800
rect 450973 328600 451477 338794
rect 450973 323200 451100 328600
rect 451400 323200 451477 328600
rect 450973 316468 451477 323200
rect 451597 336200 451857 338794
rect 451597 330800 451700 336200
rect 451800 330800 451857 336200
rect 451597 316468 451857 330800
rect 451977 336200 452499 338794
rect 451977 330800 452100 336200
rect 452400 330800 452499 336200
rect 451977 316468 452499 330800
rect 452619 328600 453767 338794
rect 452619 323200 452700 328600
rect 453700 323200 453767 328600
rect 452619 316468 453767 323200
rect 453887 336200 454617 338794
rect 453887 330800 454000 336200
rect 454500 330800 454617 336200
rect 453887 316468 454617 330800
rect 454737 328600 455241 338794
rect 454737 323200 454800 328600
rect 455100 323200 455241 328600
rect 454737 316468 455241 323200
rect 455361 336200 455621 338794
rect 455361 330800 455400 336200
rect 455500 330800 455621 336200
rect 455361 316468 455621 330800
rect 455741 336200 456263 338794
rect 455741 330800 455800 336200
rect 456200 330800 456263 336200
rect 455741 316468 456263 330800
rect 456383 328600 457531 338794
rect 456383 323200 456500 328600
rect 457500 323200 457531 328600
rect 456383 316468 457531 323200
rect 457651 336200 458381 338794
rect 457651 330800 457800 336200
rect 458300 330800 458381 336200
rect 457651 316468 458381 330800
rect 458501 328600 459005 338794
rect 458501 323200 458600 328600
rect 458900 323200 459005 328600
rect 458501 316468 459005 323200
rect 459125 336200 459385 338794
rect 459125 330800 459200 336200
rect 459300 330800 459385 336200
rect 459125 316468 459385 330800
rect 459505 336200 460027 338794
rect 459505 330800 459600 336200
rect 459900 330800 460027 336200
rect 459505 316468 460027 330800
rect 460147 328600 461295 338794
rect 460147 323200 460200 328600
rect 461200 323200 461295 328600
rect 460147 316468 461295 323200
rect 461415 336200 462145 338794
rect 461415 330800 461500 336200
rect 462000 330800 462145 336200
rect 461415 316468 462145 330800
rect 462265 328600 462769 338794
rect 462265 323200 462400 328600
rect 462700 323200 462769 328600
rect 462265 316468 462769 323200
rect 462889 336200 463149 338794
rect 462889 330800 463000 336200
rect 463100 330800 463149 336200
rect 462889 316468 463149 330800
rect 463269 336200 463791 338794
rect 463269 330800 463400 336200
rect 463700 330800 463791 336200
rect 463269 316468 463791 330800
rect 463911 328600 465059 338794
rect 463911 323200 464000 328600
rect 465000 323200 465059 328600
rect 463911 316468 465059 323200
rect 465179 336200 465909 338794
rect 465179 330800 465300 336200
rect 465800 330800 465909 336200
rect 465179 316468 465909 330800
rect 466029 328600 466533 338794
rect 466029 323200 466100 328600
rect 466400 323200 466533 328600
rect 466029 316468 466533 323200
rect 466733 336200 467653 338794
rect 466733 330800 466800 336200
rect 467600 330800 467653 336200
rect 466733 316468 467653 330800
rect 467781 328600 468681 338794
rect 467781 323200 467900 328600
rect 468600 323200 468681 328600
rect 467781 316468 468681 323200
rect 52542 315756 54180 315882
rect 37548 315630 38808 315756
rect 37548 314874 37674 315630
rect 38682 314874 38808 315630
rect 37548 314748 38808 314874
rect 52542 315504 52668 315756
rect 54054 315504 54180 315756
rect 33750 314285 49026 314545
rect 32550 308767 32810 308849
rect 32550 198350 32810 308528
rect 33150 308296 33410 308356
rect 33150 223279 33410 308123
rect 33750 257276 34010 314285
rect 34350 313811 41985 314071
rect 33695 257206 34047 257276
rect 33695 254062 33739 257206
rect 33994 254062 34047 257206
rect 33695 254010 34047 254062
rect 33126 223223 33425 223279
rect 33126 219357 33176 223223
rect 33382 219357 33425 223223
rect 33126 219314 33425 219357
rect 33150 219293 33410 219314
rect 32550 123691 32810 198151
rect 33750 199085 34010 254010
rect 34350 240476 34610 313811
rect 35028 313488 36036 313614
rect 35028 312984 35154 313488
rect 35910 312984 36036 313488
rect 35028 312858 36036 312984
rect 38386 313604 38625 313631
rect 38386 313329 38413 313604
rect 38578 313329 38625 313604
rect 41725 313623 41985 313811
rect 41725 313357 41744 313623
rect 41962 313357 41985 313623
rect 41725 313337 41985 313357
rect 42714 313614 43344 313740
rect 38386 308767 38625 313329
rect 42714 312858 42840 313614
rect 43218 312858 43344 313614
rect 42714 312732 43344 312858
rect 43974 313687 44478 313740
rect 43974 313428 44030 313687
rect 44407 313428 44478 313687
rect 43974 313362 44478 313428
rect 45418 313601 45657 313668
rect 48766 313649 49026 314285
rect 43974 311220 44226 313362
rect 45418 313339 45467 313601
rect 45631 313339 45657 313601
rect 48764 313634 49026 313649
rect 48764 313364 48779 313634
rect 49011 313364 49026 313634
rect 52542 314496 54180 315504
rect 63630 315630 65142 315756
rect 63630 315378 63756 315630
rect 65016 315378 65142 315630
rect 52542 313740 52668 314496
rect 54054 313740 54180 314496
rect 52542 313614 54180 313740
rect 58464 314496 59472 314622
rect 58464 313740 58590 314496
rect 59346 313740 59472 314496
rect 58464 313614 59472 313740
rect 63630 314496 65142 315378
rect 63630 313740 63756 314496
rect 65016 313740 65142 314496
rect 63630 313614 65142 313740
rect 68544 314496 69552 314622
rect 68544 313740 68670 314496
rect 69426 313740 69552 314496
rect 48764 313345 49026 313364
rect 43974 311094 44478 311220
rect 42714 310842 43344 310968
rect 42714 310338 42840 310842
rect 43218 310338 43344 310842
rect 42714 310212 43344 310338
rect 43974 310212 44100 311094
rect 44352 310212 44478 311094
rect 43974 310086 44478 310212
rect 38386 308474 38625 308528
rect 45418 308767 45657 313339
rect 50268 312393 58126 312396
rect 50268 312160 50283 312393
rect 50882 312160 58126 312393
rect 50268 312156 58126 312160
rect 49896 310842 50526 310968
rect 49896 310338 50022 310842
rect 50400 310338 50526 310842
rect 49896 310212 50526 310338
rect 57886 310424 58126 312156
rect 57886 310206 57903 310424
rect 58105 310206 58126 310424
rect 57886 310183 58126 310206
rect 50526 309582 51408 309708
rect 50526 309078 50652 309582
rect 51282 309078 51408 309582
rect 50526 308952 51408 309078
rect 58464 309582 58968 313614
rect 60228 313362 61362 313488
rect 60228 313110 60354 313362
rect 61236 313110 61362 313362
rect 60228 311724 61362 313110
rect 60228 311472 60354 311724
rect 61236 311472 61362 311724
rect 60228 309834 61362 311472
rect 64386 312732 65520 312858
rect 64386 312480 64512 312732
rect 65394 312480 65520 312732
rect 64386 311094 65520 312480
rect 64386 310842 64512 311094
rect 65394 310842 65520 311094
rect 68544 311220 69552 313740
rect 68544 310968 68670 311220
rect 69426 310968 69552 311220
rect 68544 310842 69552 310968
rect 64386 310212 64512 310716
rect 65394 310212 65520 310716
rect 64386 310086 65520 310212
rect 58464 308952 58590 309582
rect 58842 308952 58968 309582
rect 58464 308826 58968 308952
rect 59220 309582 61488 309834
rect 59220 308826 59346 309582
rect 61362 308826 61488 309582
rect 45418 308514 45657 308528
rect 59220 307692 61488 308826
rect 59220 307062 59346 307692
rect 61362 307062 61488 307692
rect 59220 306936 61488 307062
rect 57834 288162 60480 288288
rect 57834 287910 57960 288162
rect 60354 287910 60480 288162
rect 54810 286272 55944 286398
rect 54810 285642 54936 286272
rect 55818 285642 55944 286272
rect 49140 284886 50274 285012
rect 49140 284256 49266 284886
rect 50148 284256 50274 284886
rect 49140 283951 50274 284256
rect 49140 283673 49186 283951
rect 50234 283673 50274 283951
rect 49140 283626 50274 283673
rect 54810 283944 55944 285642
rect 57834 286272 60480 287910
rect 57834 285642 57960 286272
rect 60354 285642 60480 286272
rect 57834 285516 60480 285642
rect 54810 283680 54858 283944
rect 55884 283680 55944 283944
rect 54810 283626 55944 283680
rect 34950 282082 35210 282159
rect 34295 240406 34647 240476
rect 34295 237262 34339 240406
rect 34594 237262 34647 240406
rect 34295 237210 34647 237262
rect 34950 237882 35210 281649
rect 34950 206876 35210 237449
rect 35550 249475 35810 249671
rect 34895 206806 35247 206876
rect 34895 203662 34939 206806
rect 35194 203662 35247 206806
rect 34895 203610 35247 203662
rect 35550 205875 35810 248888
rect 58464 247968 59346 248094
rect 58464 247086 58590 247968
rect 59220 247086 59346 247968
rect 58464 246960 59346 247086
rect 60102 246330 60982 246456
rect 60102 245448 60228 246330
rect 60858 245448 60982 246330
rect 60102 245322 60982 245448
rect 63756 244692 64764 244818
rect 63756 243936 63882 244692
rect 64638 243936 64764 244692
rect 63756 243882 64764 243936
rect 44334 243288 44526 243326
rect 44334 242122 44526 242190
rect 67158 243180 68040 243306
rect 67158 242298 67284 243180
rect 67914 242298 68040 243180
rect 67158 242172 68040 242298
rect 65638 241794 67024 241920
rect 65638 241290 65764 241794
rect 66898 241290 67024 241794
rect 65638 241164 67024 241290
rect 33750 124240 34010 198886
rect 34950 195219 35198 203610
rect 34950 195082 35210 195219
rect 34950 194522 35210 194649
rect 35550 190076 35810 205288
rect 36750 240127 65108 240387
rect 36150 197670 36410 197740
rect 35495 190006 35847 190076
rect 35495 186862 35539 190006
rect 35794 186862 35847 190006
rect 35495 186810 35847 186862
rect 35550 163075 35810 186810
rect 36150 173276 36410 197377
rect 36095 173206 36447 173276
rect 36095 170062 36139 173206
rect 36394 170062 36447 173206
rect 36095 170010 36447 170062
rect 35550 162239 35810 162488
rect 36750 156476 37010 240127
rect 49644 239904 51786 240030
rect 49644 239778 49770 239904
rect 51660 239778 51786 239904
rect 49644 239652 51786 239778
rect 64848 239346 65108 240127
rect 64848 238630 64857 239346
rect 65097 238630 65108 239346
rect 64848 238597 65108 238630
rect 66276 233604 66780 233730
rect 66276 232596 66402 233604
rect 66654 232596 66780 233604
rect 66276 232470 66780 232596
rect 72324 229320 73710 229446
rect 72324 228690 72450 229320
rect 73584 228690 73710 229320
rect 72324 228564 73710 228690
rect 65268 226674 66654 226800
rect 65268 225792 65394 226674
rect 66528 225792 66654 226674
rect 65268 225666 66654 225792
rect 72828 209538 73710 209664
rect 72828 208656 72954 209538
rect 73584 208656 73710 209538
rect 72828 208530 73710 208656
rect 79254 207942 79758 208026
rect 79254 206980 79331 207942
rect 79685 206980 79758 207942
rect 79254 206892 79758 206980
rect 74306 205722 74654 205762
rect 74306 205038 74345 205722
rect 74614 205038 74654 205722
rect 74306 204996 74654 205038
rect 73080 200970 87696 201096
rect 73080 199710 73206 200970
rect 73710 200466 82404 200970
rect 73710 199710 73836 200466
rect 82278 200340 82404 200466
rect 87570 200340 87696 200970
rect 82278 200214 87696 200340
rect 73080 199584 73836 199710
rect 70686 198850 71442 198976
rect 70686 198094 70812 198850
rect 71316 198094 71442 198850
rect 70686 197968 71442 198094
rect 49789 197117 51889 197164
rect 49789 196869 49829 197117
rect 51830 196869 51889 197117
rect 49789 196826 51889 196869
rect 68922 193032 69678 193158
rect 68922 192402 69048 193032
rect 69552 192402 69678 193032
rect 68922 192276 69678 192402
rect 66024 190008 66906 190134
rect 66024 189252 66150 190008
rect 66780 189252 66906 190008
rect 66024 189126 66906 189252
rect 65646 184212 67032 184338
rect 65646 183078 65772 184212
rect 66906 183078 67032 184212
rect 65646 182952 67032 183078
rect 73206 167202 79758 167328
rect 73206 166446 73332 167202
rect 74088 166446 74970 167202
rect 79632 166446 79758 167202
rect 73206 166320 79758 166446
rect 79380 165312 80010 165438
rect 79380 164178 79506 165312
rect 79884 164178 80010 165312
rect 79380 164052 80010 164178
rect 80766 162036 81648 162288
rect 80766 161532 80892 162036
rect 81522 161532 81648 162036
rect 70878 156752 71846 156878
rect 70878 156500 70964 156752
rect 71720 156500 71846 156752
rect 36695 156406 37047 156476
rect 36695 153262 36739 156406
rect 36994 153262 37047 156406
rect 70878 156374 71846 156500
rect 71986 156744 72954 156870
rect 71986 156492 72072 156744
rect 72828 156492 72954 156744
rect 71986 156366 72954 156492
rect 80766 154980 81648 161532
rect 80766 154224 80892 154980
rect 81522 154224 81648 154980
rect 80766 154098 81648 154224
rect 36695 153210 37047 153262
rect 51282 153468 52920 153594
rect 51282 152838 51408 153468
rect 52794 153342 83158 153468
rect 52794 152964 70938 153342
rect 73710 152964 83158 153342
rect 52794 152838 83158 152964
rect 51282 152712 52920 152838
rect 59724 151956 60354 152082
rect 59724 149562 59850 151956
rect 60228 149562 60354 151956
rect 59724 149436 60354 149562
rect 59850 130536 60102 149436
rect 81144 146412 81774 146538
rect 81144 142380 81270 146412
rect 81648 142380 81774 146412
rect 82528 145040 83158 152838
rect 321000 149736 321600 149836
rect 321000 149336 321100 149736
rect 321500 149336 321600 149736
rect 321000 149236 321600 149336
rect 321000 148736 321600 148836
rect 321000 148336 321100 148736
rect 321500 148336 321600 148736
rect 321000 148236 321600 148336
rect 82432 144978 83216 145040
rect 82432 144633 82494 144978
rect 83152 144633 83216 144978
rect 82432 144592 83216 144633
rect 81144 142254 81774 142380
rect 89152 139328 90832 139440
rect 89152 138432 89264 139328
rect 90720 138432 90832 139328
rect 89152 138320 90832 138432
rect 60858 135828 61488 135954
rect 60858 133560 60984 135828
rect 61362 133560 61488 135828
rect 60858 133434 61488 133560
rect 275800 133700 276600 133800
rect 275800 133100 275900 133700
rect 276500 133100 276600 133700
rect 275800 133000 276600 133100
rect 72188 132804 73196 132930
rect 72188 132174 72314 132804
rect 73070 132174 73196 132804
rect 62622 131292 65772 131418
rect 62622 131040 62748 131292
rect 65646 131040 65772 131292
rect 62622 130914 65772 131040
rect 72188 130536 73196 132174
rect 121464 132426 206136 132552
rect 121464 131040 202860 132426
rect 74592 130662 80136 130788
rect 74592 130536 74718 130662
rect 59850 130511 61992 130536
rect 59850 130057 59875 130511
rect 60078 130477 61992 130511
rect 60078 130057 61634 130477
rect 59850 130051 61634 130057
rect 61874 130051 61992 130477
rect 59850 130032 61992 130051
rect 62622 130410 74718 130536
rect 62622 130158 62748 130410
rect 65646 130158 74718 130410
rect 62622 130032 74718 130158
rect 80010 130032 80136 130662
rect 59850 127764 60102 130032
rect 74592 129906 80136 130032
rect 121464 130032 121590 131040
rect 124866 130032 202860 131040
rect 206010 130032 206136 132426
rect 275800 132300 276600 132400
rect 275800 131700 275900 132300
rect 276500 131700 276600 132300
rect 275800 131600 276600 131700
rect 121464 129906 206136 130032
rect 59724 127638 60228 127764
rect 59724 127386 59850 127638
rect 60102 127386 60228 127638
rect 59724 127260 60228 127386
rect 60984 127008 61992 127134
rect 60984 126630 61110 127008
rect 61866 126630 61992 127008
rect 60984 126504 61992 126630
rect 33750 123980 37300 124240
rect 32550 123431 36688 123691
rect 34524 116046 35532 116172
rect 34524 114912 34650 116046
rect 35406 114912 35532 116046
rect 34524 114786 35532 114912
rect 36288 71921 36688 123431
rect 37040 110632 37300 123980
rect 98784 111888 102816 112014
rect 74466 111636 80136 111762
rect 37040 110609 73710 110632
rect 37040 110390 73470 110609
rect 73693 110390 73710 110609
rect 37040 110372 73710 110390
rect 74466 110502 74592 111636
rect 80010 111006 80136 111636
rect 80010 110880 90972 111006
rect 80010 110502 90468 110880
rect 90846 110502 90972 110880
rect 74466 110376 90972 110502
rect 98784 109746 98910 111888
rect 37548 109620 98910 109746
rect 37548 108612 37674 109620
rect 38556 109116 91476 109620
rect 38556 108738 66906 109116
rect 67536 108738 91476 109116
rect 91728 108738 98910 109620
rect 38556 108612 98910 108738
rect 102690 108612 102816 111888
rect 37548 108486 102816 108612
rect 103950 110376 114282 110502
rect 103950 107982 104076 110376
rect 38304 107856 104076 107982
rect 38304 107604 74340 107856
rect 38304 107352 65898 107604
rect 38304 106974 59598 107352
rect 60606 107226 65898 107352
rect 66528 107352 74340 107604
rect 75096 107352 92484 107856
rect 92988 107352 104076 107856
rect 66528 107226 104076 107352
rect 60606 107100 104076 107226
rect 107730 107100 108864 110376
rect 114156 107100 114282 110376
rect 60606 106974 114282 107100
rect 38304 106722 107856 106974
rect 98784 84879 104328 85005
rect 98784 82782 98910 84879
rect 104202 82782 104328 84879
rect 98784 82656 104328 82782
rect 477200 79400 477800 79500
rect 477200 79000 477300 79400
rect 477700 79000 477800 79400
rect 477200 78900 477800 79000
rect 477200 78400 477800 78500
rect 477200 78000 477300 78400
rect 477700 78000 477800 78400
rect 477200 77900 477800 78000
rect 472400 75600 478000 75800
rect 135946 72828 140986 72954
rect 113148 72072 114030 72198
rect 36288 71868 36848 71921
rect 36288 71511 36848 71588
rect 113148 71442 113274 72072
rect 113904 71442 114030 72072
rect 113148 71316 114030 71442
rect 135946 71442 136072 72828
rect 140860 71442 140986 72828
rect 135946 71316 140986 71442
rect 96894 70938 106344 71064
rect 96894 69426 97020 70938
rect 106218 69426 106344 70938
rect 96894 69300 106344 69426
rect 211176 61614 213192 61740
rect 211176 59220 211302 61614
rect 213066 59220 213192 61614
rect 268380 61362 283248 61488
rect 268380 59472 268506 61362
rect 283122 59472 283248 61362
rect 472400 61200 472600 75600
rect 477800 61200 478000 75600
rect 472400 61000 478000 61200
rect 268380 59346 283248 59472
rect 211176 58022 213192 59220
rect 285200 58600 300000 58800
rect 34400 57600 36400 57800
rect 34400 43200 34600 57600
rect 36200 43200 36400 57600
rect 211176 55766 215192 58022
rect 199000 53800 204646 54000
rect 199000 51600 199200 53800
rect 204464 51600 204646 53800
rect 199000 51400 204646 51600
rect 205266 53800 211000 54000
rect 205266 51600 205440 53800
rect 210800 51600 211000 53800
rect 205266 51400 211000 51600
rect 96138 50526 107604 50652
rect 96138 47754 96264 50526
rect 107478 47754 107604 50526
rect 96138 47628 107604 47754
rect 34400 43000 36400 43200
rect 213176 41832 215192 55766
rect 285200 53400 285400 58600
rect 299800 53400 300000 58600
rect 285200 53200 300000 53400
rect 317800 52300 318600 52400
rect 317800 51700 317900 52300
rect 318500 51700 318600 52300
rect 317800 51600 318600 51700
rect 317800 51100 318600 51200
rect 317800 50500 317900 51100
rect 318500 50500 318600 51100
rect 317800 50400 318600 50500
rect 480400 45100 481200 45200
rect 480400 44500 480500 45100
rect 481100 44500 481200 45100
rect 480400 44400 481200 44500
rect 480400 43700 481200 43800
rect 480400 43100 480500 43700
rect 481100 43100 481200 43700
rect 480400 43000 481200 43100
rect 231600 42200 246400 42400
rect 231600 41832 231800 42200
rect 59700 41700 60500 41800
rect 59700 41100 59800 41700
rect 60400 41100 60500 41700
rect 59700 41000 60500 41100
rect 59700 40500 60500 40600
rect 59700 39900 59800 40500
rect 60400 39900 60500 40500
rect 59700 39800 60500 39900
rect 213176 39816 231800 41832
rect 231600 37200 231800 39816
rect 246200 37200 246400 42200
rect 231600 37000 246400 37200
rect 102200 35400 117000 35600
rect 102200 33800 102400 35400
rect 116800 33800 117000 35400
rect 102200 33600 117000 33800
<< viatp >>
rect 33600 366000 34600 380400
rect 332154 380250 332744 380778
rect 427400 374200 441800 375800
rect 444200 374200 447000 375800
rect 452600 374200 458600 375800
rect 467000 374200 481400 375800
rect 41076 366786 44604 368424
rect 33600 349200 34600 363600
rect 60102 366786 62748 368046
rect 63504 366912 64764 367542
rect 320796 365354 322407 365486
rect 320796 364604 322686 365354
rect 328600 364800 329200 365400
rect 328600 363400 329200 364000
rect 322056 361872 323316 362502
rect 63126 358092 63378 358470
rect 66150 360360 66780 361620
rect 326340 361242 329364 362880
rect 65394 357714 65646 358470
rect 334600 360800 346000 362200
rect 470300 373000 470800 373500
rect 471500 373000 472000 373500
rect 472600 349200 477800 363600
rect 37800 335916 40068 336798
rect 49518 335916 51786 336798
rect 61992 335916 64260 336798
rect 328200 323200 329000 328600
rect 329300 330800 329900 336200
rect 330200 323200 330300 328600
rect 330600 330800 330700 336200
rect 331000 330800 331300 336200
rect 331600 323200 332600 328600
rect 332900 330800 333400 336200
rect 333700 323200 334000 328600
rect 334300 330800 334400 336200
rect 334700 330800 335000 336200
rect 335400 323200 336400 328600
rect 336700 330800 337200 336200
rect 337500 323200 337800 328600
rect 338100 330800 338200 336200
rect 338500 330800 338800 336200
rect 339200 323200 340200 328600
rect 340500 330800 341000 336200
rect 341300 323200 341600 328600
rect 341900 330800 342000 336200
rect 342300 330800 342600 336200
rect 342900 323200 343900 328600
rect 344200 330800 344700 336200
rect 345000 323200 345300 328600
rect 345600 330800 345700 336200
rect 346100 330800 346400 336200
rect 346700 323200 347700 328600
rect 348000 330800 348500 336200
rect 348800 323200 349100 328600
rect 349400 330800 349500 336200
rect 349800 330800 350100 336200
rect 350400 323200 351400 328600
rect 351700 330800 352200 336200
rect 352600 323200 352900 328600
rect 353200 330800 353300 336200
rect 353600 330800 353900 336200
rect 354200 323200 355200 328600
rect 355500 330800 356000 336200
rect 356300 323200 356600 328600
rect 356900 330800 357000 336200
rect 357300 330800 357600 336200
rect 358000 323200 359000 328600
rect 359300 330800 359800 336200
rect 360100 323200 360400 328600
rect 360700 330800 360800 336200
rect 361100 330800 361400 336200
rect 361700 323200 362700 328600
rect 363000 330800 363500 336200
rect 363900 323200 364200 328600
rect 364500 330800 364600 336200
rect 364900 330800 365200 336200
rect 365500 323200 366500 328600
rect 366800 330800 367300 336200
rect 367600 323200 367900 328600
rect 368200 330800 368300 336200
rect 368600 330800 368900 336200
rect 369200 323200 370200 328600
rect 370600 330800 371100 336200
rect 371400 323200 371700 328600
rect 372000 330800 372100 336200
rect 372400 330800 372700 336200
rect 373000 323200 374000 328600
rect 374300 330800 374800 336200
rect 375100 323200 375400 328600
rect 375800 330800 375900 336200
rect 376200 330800 376500 336200
rect 376800 323200 377800 328600
rect 378100 330800 378600 336200
rect 378900 323200 379200 328600
rect 379500 330800 379600 336200
rect 379900 330800 380200 336200
rect 380600 323200 381600 328600
rect 381800 330800 382300 336200
rect 382700 323200 383000 328600
rect 383300 330800 383400 336200
rect 383700 330800 384000 336200
rect 384300 323200 385300 328600
rect 385600 330800 386100 336200
rect 386400 323200 386700 328600
rect 387100 330800 387200 336200
rect 387500 330800 387800 336200
rect 388100 323200 389100 328600
rect 389400 330800 389900 336200
rect 390200 323200 390500 328600
rect 390800 330800 391000 336200
rect 391300 323200 391700 328600
rect 392200 330800 392500 336200
rect 392800 323200 393800 328600
rect 394300 330800 395800 336200
rect 396100 323200 396400 328600
rect 396800 330800 397800 336200
rect 398200 323200 400000 328600
rect 400600 330800 401800 336200
rect 402300 323200 403300 328600
rect 403600 323200 404600 328600
rect 404900 330800 405400 336200
rect 405700 323200 406200 328600
rect 406500 330800 406600 336200
rect 406900 330800 407300 336200
rect 407500 323200 408500 328600
rect 408800 330800 409300 336200
rect 409700 323200 410000 328600
rect 410300 330800 410400 336200
rect 410700 330800 411000 336200
rect 411300 323200 412300 328600
rect 412600 330800 413100 336200
rect 413400 323200 413700 328600
rect 414000 330800 414100 336200
rect 414400 330800 414700 336200
rect 415100 323200 416100 328600
rect 416400 330800 416900 336200
rect 417200 323200 417500 328600
rect 417800 330800 417900 336200
rect 418200 330800 418500 336200
rect 418800 323200 419800 328600
rect 420100 330800 420600 336200
rect 420900 323200 421200 328600
rect 421600 330800 421700 336200
rect 422000 330800 422300 336200
rect 422600 323200 423600 328600
rect 423900 330800 424400 336200
rect 424700 323200 425000 328600
rect 425300 330800 425400 336200
rect 425700 330800 426000 336200
rect 426400 323200 427400 328600
rect 427600 330800 428100 336200
rect 428500 323200 428800 328600
rect 429100 330800 429200 336200
rect 429500 330800 429800 336200
rect 430100 323200 431100 328600
rect 431400 330800 431900 336200
rect 432300 323200 432600 328600
rect 432800 330800 432900 336200
rect 433300 330800 433600 336200
rect 433900 323200 434900 328600
rect 435200 330800 435700 336200
rect 436000 323200 436300 328600
rect 436600 330800 436700 336200
rect 437000 330800 437300 336200
rect 437600 323200 438600 328600
rect 438900 330800 439400 336200
rect 439800 323200 440100 328600
rect 440400 330800 440500 336200
rect 440800 330800 441100 336200
rect 441400 323200 442400 328600
rect 442700 330800 443200 336200
rect 443500 323200 443800 328600
rect 444100 330800 444200 336200
rect 444600 330800 444900 336200
rect 445200 323200 446200 328600
rect 446500 330800 447000 336200
rect 447300 323200 447600 328600
rect 447900 330800 448000 336200
rect 448300 330800 448600 336200
rect 448900 323200 449900 328600
rect 450200 330800 450700 336200
rect 451100 323200 451400 328600
rect 451700 330800 451800 336200
rect 452100 330800 452400 336200
rect 452700 323200 453700 328600
rect 454000 330800 454500 336200
rect 454800 323200 455100 328600
rect 455400 330800 455500 336200
rect 455800 330800 456200 336200
rect 456500 323200 457500 328600
rect 457800 330800 458300 336200
rect 458600 323200 458900 328600
rect 459200 330800 459300 336200
rect 459600 330800 459900 336200
rect 460200 323200 461200 328600
rect 461500 330800 462000 336200
rect 462400 323200 462700 328600
rect 463000 330800 463100 336200
rect 463400 330800 463700 336200
rect 464000 323200 465000 328600
rect 465300 330800 465800 336200
rect 466100 323200 466400 328600
rect 466800 330800 467600 336200
rect 467900 323200 468600 328600
rect 37674 315378 38682 315630
rect 37674 314874 38682 315378
rect 35154 312984 35910 313488
rect 42840 312858 43218 313614
rect 52668 313740 54054 314496
rect 58590 313740 59346 314496
rect 63756 313740 65016 314496
rect 68670 313740 69426 314496
rect 42840 310338 43218 310842
rect 44100 310212 44352 311094
rect 50022 310338 50400 310842
rect 50652 309078 51282 309582
rect 64512 310842 65394 311094
rect 64512 310716 65394 310842
rect 64512 310212 65394 310716
rect 59346 308826 61362 309582
rect 54936 285642 55818 286272
rect 49266 284256 50148 284886
rect 57960 285642 60354 286272
rect 58590 247086 59220 247968
rect 60228 245448 60858 246330
rect 63882 243936 64638 244692
rect 44334 242190 44526 243288
rect 67284 242298 67914 243180
rect 65764 241290 66898 241794
rect 49770 239778 51660 239904
rect 66402 232596 66654 233604
rect 72450 228690 73584 229320
rect 65394 225792 66528 226674
rect 72954 208656 73584 209538
rect 79331 206980 79685 207942
rect 74345 205038 74614 205722
rect 82404 200340 87570 200970
rect 70812 198094 71316 198850
rect 49829 196869 51830 197117
rect 69048 192402 69552 193032
rect 66150 189252 66780 190008
rect 65772 183078 66906 184212
rect 74970 166446 79632 167202
rect 79506 164178 79884 165312
rect 70964 156500 71720 156752
rect 72072 156492 72828 156744
rect 80892 154224 81522 154980
rect 70938 152964 73710 153342
rect 59850 149562 60228 151956
rect 81270 142380 81648 146412
rect 321100 149336 321500 149736
rect 321100 148336 321500 148736
rect 89264 138432 90720 139328
rect 60984 133560 61362 135828
rect 275900 133100 276500 133700
rect 62748 131040 65646 131292
rect 74718 130032 80010 130662
rect 121590 130032 124866 131040
rect 202860 130032 206010 132426
rect 275900 131700 276500 132300
rect 61110 126630 61866 127008
rect 34650 114912 35406 116046
rect 74592 110502 80010 111636
rect 98910 108612 102690 111888
rect 108864 107100 114156 110376
rect 98910 82782 99920 84879
rect 99920 82782 100344 84879
rect 100344 82782 101224 84879
rect 101224 82782 101680 84879
rect 101680 82782 102540 84879
rect 102540 82782 102967 84879
rect 102967 82782 104202 84879
rect 477300 79000 477700 79400
rect 477300 78000 477700 78400
rect 113274 71442 113904 72072
rect 136072 71442 140860 72828
rect 97020 69426 106218 70938
rect 211302 59220 213066 61614
rect 268506 59472 283122 61362
rect 472600 61200 477800 75600
rect 34600 43200 36200 57600
rect 199200 51600 204464 53800
rect 205440 51600 210800 53800
rect 96264 47754 97476 50526
rect 97476 47754 97964 50526
rect 97964 47754 99320 50526
rect 99320 47754 99742 50526
rect 99742 47754 100567 50526
rect 100567 47754 100966 50526
rect 100966 47754 101841 50526
rect 101841 47754 102284 50526
rect 102284 47754 103006 50526
rect 103006 47754 103453 50526
rect 103453 47754 104649 50526
rect 104649 47754 105096 50526
rect 105096 47754 105822 50526
rect 105822 47754 106276 50526
rect 106276 47754 107478 50526
rect 285400 53400 299800 58600
rect 317900 51700 318500 52300
rect 317900 50500 318500 51100
rect 480500 44500 481100 45100
rect 480500 43100 481100 43700
rect 59800 41100 60400 41700
rect 59800 39900 60400 40500
rect 231800 37200 246200 42200
rect 102400 33800 116800 35400
<< metaltp >>
rect 332100 380778 332806 380830
rect 82256 380634 331280 380694
rect 33400 380400 34800 380600
rect 33400 366000 33600 380400
rect 34600 372331 34800 380400
rect 82256 379520 319364 380634
rect 324824 379520 331280 380634
rect 332100 380250 332154 380778
rect 332744 380250 332806 380778
rect 332100 380188 332806 380250
rect 82256 379448 331280 379520
rect 84217 379018 84356 379448
rect 88747 379018 88886 379448
rect 93277 379018 93416 379448
rect 97807 379018 97946 379448
rect 102337 379018 102476 379448
rect 106867 379018 107006 379448
rect 111397 379018 111536 379448
rect 115927 379018 116066 379448
rect 120457 379018 120596 379448
rect 124987 379018 125126 379448
rect 129517 379018 129656 379448
rect 134047 379018 134186 379448
rect 138577 379018 138716 379448
rect 143107 379018 143246 379448
rect 147637 379018 147776 379448
rect 152167 379018 152306 379448
rect 156697 379018 156836 379448
rect 161227 379018 161366 379448
rect 165757 379018 165896 379448
rect 170287 379018 170426 379448
rect 174817 379018 174956 379448
rect 179347 379018 179486 379448
rect 183877 379018 184016 379448
rect 188407 379018 188546 379448
rect 192937 379018 193076 379448
rect 197467 379018 197606 379448
rect 201997 379018 202136 379448
rect 206527 379018 206666 379448
rect 211057 379018 211196 379448
rect 215587 379018 215726 379448
rect 220117 379018 220256 379448
rect 224647 379018 224786 379448
rect 229177 379018 229316 379448
rect 233707 379018 233846 379448
rect 238237 379018 238376 379448
rect 242767 379018 242906 379448
rect 247297 379018 247436 379448
rect 251827 379018 251966 379448
rect 256357 379018 256496 379448
rect 260887 379018 261026 379448
rect 265417 379018 265556 379448
rect 269947 379018 270086 379448
rect 274477 379018 274616 379448
rect 279007 379018 279146 379448
rect 283537 379018 283676 379448
rect 288067 379018 288206 379448
rect 292597 379018 292736 379448
rect 297127 379018 297266 379448
rect 301657 379018 301796 379448
rect 306187 379018 306326 379448
rect 310717 379018 310856 379448
rect 315247 379018 315386 379448
rect 319777 379018 319916 379448
rect 324307 379018 324446 379448
rect 328837 379018 328976 379448
rect 34600 368424 74544 372331
rect 34600 366786 41076 368424
rect 44604 368046 74544 368424
rect 44604 366786 60102 368046
rect 62748 367542 74544 368046
rect 62748 366912 63504 367542
rect 64764 366912 74544 367542
rect 62748 366786 74544 366912
rect 34600 366731 74544 366786
rect 80144 366731 80811 372331
rect 34600 366000 34800 366731
rect 33400 365800 34800 366000
rect 86437 364731 86577 366088
rect 90967 364731 91107 366088
rect 95497 364731 95637 366088
rect 100027 364731 100167 366088
rect 104557 364731 104697 366088
rect 109087 364731 109227 366152
rect 113617 364731 113757 366152
rect 118147 364731 118287 366152
rect 122677 364731 122817 366152
rect 127207 364731 127347 366152
rect 131737 364731 131877 366152
rect 136267 364731 136407 366152
rect 140797 364731 140937 366152
rect 145327 364731 145467 366152
rect 149857 364731 149997 366152
rect 154387 364731 154527 366152
rect 158917 364731 159057 366152
rect 163447 364731 163587 366152
rect 167977 364731 168117 366152
rect 172507 364731 172647 366152
rect 177037 364731 177177 366152
rect 181567 364731 181707 366152
rect 186097 364731 186237 366152
rect 190627 364731 190767 366152
rect 195157 364731 195297 366152
rect 199687 364731 199827 366152
rect 204217 364731 204357 366152
rect 208747 364731 208887 366152
rect 213277 364731 213417 366152
rect 217807 364731 217947 366152
rect 222337 364731 222477 366152
rect 226867 364731 227007 366152
rect 231397 364731 231537 366152
rect 235927 364731 236067 366152
rect 240457 364731 240597 366152
rect 244987 364731 245127 366152
rect 249517 364731 249657 366152
rect 254047 364731 254187 366152
rect 258577 364731 258717 366152
rect 263107 364731 263247 366152
rect 267637 364731 267777 366152
rect 272167 364731 272307 366152
rect 276697 364731 276837 366152
rect 281227 364731 281367 366152
rect 285757 364731 285897 366152
rect 290287 364731 290427 366152
rect 294817 364731 294957 366152
rect 299347 364731 299487 366152
rect 303877 364731 304017 366152
rect 308407 364731 308547 366152
rect 312937 364731 313077 366152
rect 317467 364731 317607 366152
rect 321997 365981 322137 366080
rect 321997 365841 323251 365981
rect 320670 365486 322812 365612
rect 33400 363600 82144 364731
rect 33400 349200 33600 363600
rect 34600 361620 82144 363600
rect 34600 360360 66150 361620
rect 66780 360360 82144 361620
rect 34600 359131 82144 360360
rect 87744 359131 108864 364731
rect 109620 359131 128772 364731
rect 129528 359131 148680 364731
rect 149436 359131 168588 364731
rect 169344 359131 188496 364731
rect 189252 359131 208404 364731
rect 209160 359131 228312 364731
rect 229068 359131 248220 364731
rect 248976 359131 268128 364731
rect 268884 359131 288036 364731
rect 288792 364072 319018 364731
rect 320670 364604 320796 365486
rect 322686 364604 322812 365486
rect 320670 364486 322812 364604
rect 323111 364084 323251 365841
rect 326527 364084 326667 366152
rect 328837 365500 328977 366100
rect 328500 365400 329300 365500
rect 328500 364800 328600 365400
rect 329200 364800 329300 365400
rect 328500 364700 329300 364800
rect 328500 364084 329300 364100
rect 331057 364084 331197 366152
rect 332180 364084 332703 380188
rect 447006 379208 452606 379484
rect 447006 376000 447210 379208
rect 427200 375800 442000 376000
rect 427200 374200 427400 375800
rect 441800 374200 442000 375800
rect 427200 374000 442000 374200
rect 444000 375800 447210 376000
rect 444000 374200 444200 375800
rect 447000 374222 447210 375800
rect 452272 376000 452606 379208
rect 452272 375800 458800 376000
rect 452272 374222 452600 375800
rect 447000 374200 452600 374222
rect 458600 374200 458800 375800
rect 444000 374004 458800 374200
rect 444000 374000 447122 374004
rect 452600 374000 458800 374004
rect 466800 375800 481600 376000
rect 466800 374200 467000 375800
rect 481400 374200 481600 375800
rect 466800 374000 481600 374200
rect 432915 373543 436452 374000
rect 467550 373543 469232 374000
rect 470200 373543 470900 373600
rect 419137 373500 470900 373543
rect 419137 373031 470300 373500
rect 419447 372638 419587 373031
rect 423977 372638 424117 373031
rect 428507 372638 428647 373031
rect 433037 372638 433177 373031
rect 437567 372638 437707 373031
rect 442097 372638 442237 373031
rect 446627 372638 446767 373031
rect 451157 372638 451297 373031
rect 455687 372638 455827 373031
rect 460217 372638 460357 373031
rect 464747 372638 464887 373031
rect 469277 372638 469417 373031
rect 470200 373000 470300 373031
rect 470800 373000 470900 373500
rect 470200 372900 470900 373000
rect 471400 373500 472100 373600
rect 471400 373000 471500 373500
rect 472000 373000 472100 373500
rect 471400 372900 472100 373000
rect 471497 372600 471637 372900
rect 323111 364072 332703 364084
rect 288792 364000 332703 364072
rect 288792 363400 328600 364000
rect 329200 363400 332703 364000
rect 288792 362938 332703 363400
rect 472400 363600 478000 363800
rect 288792 362880 329490 362938
rect 288792 362502 326340 362880
rect 288792 361872 322056 362502
rect 323316 361872 326340 362502
rect 288792 361242 326340 361872
rect 329364 361242 329490 362880
rect 288792 361116 329490 361242
rect 334400 362200 346200 362400
rect 288792 359131 325000 361116
rect 334400 360800 334600 362200
rect 346000 360800 346200 362200
rect 334400 360600 346200 360800
rect 34600 349200 34800 359131
rect 35658 358470 73962 358596
rect 35658 357588 35784 358470
rect 37170 358092 63126 358470
rect 63378 358092 65394 358470
rect 37170 357714 65394 358092
rect 65646 357714 73962 358470
rect 37170 357588 73962 357714
rect 35658 357462 73962 357588
rect 33400 349000 34800 349200
rect 37044 336798 87696 336924
rect 37044 335916 37800 336798
rect 40068 335916 49518 336798
rect 51786 335916 61992 336798
rect 64260 335916 82278 336798
rect 87570 335916 87696 336798
rect 37044 335790 87696 335916
rect 316853 336342 317988 336344
rect 319400 336342 325000 359131
rect 472400 349200 472600 363600
rect 477800 349200 478000 363600
rect 472400 349000 478000 349200
rect 421667 336342 421807 342429
rect 426197 336342 426337 342490
rect 430727 336342 430867 342429
rect 435257 336342 435397 342429
rect 439787 336342 439927 342429
rect 444317 336342 444457 342429
rect 448847 336342 448987 342429
rect 453377 336342 453517 342429
rect 457907 336342 458047 342429
rect 462437 336342 462577 342429
rect 466967 336342 467107 342429
rect 471497 336342 471637 342429
rect 316853 336200 447000 336342
rect 452600 336200 472387 336342
rect 316853 330800 329300 336200
rect 329900 330800 330600 336200
rect 330700 330800 331000 336200
rect 331300 330800 332900 336200
rect 333400 330800 334300 336200
rect 334400 330800 334700 336200
rect 335000 330800 336700 336200
rect 337200 330800 338100 336200
rect 338200 330800 338500 336200
rect 338800 330800 340500 336200
rect 341000 330800 341900 336200
rect 342000 330800 342300 336200
rect 342600 330800 344200 336200
rect 344700 330800 345600 336200
rect 345700 330800 346100 336200
rect 346400 330800 348000 336200
rect 348500 330800 349400 336200
rect 349500 330800 349800 336200
rect 350100 330800 351700 336200
rect 352200 330800 353200 336200
rect 353300 330800 353600 336200
rect 353900 330800 355500 336200
rect 356000 330800 356900 336200
rect 357000 330800 357300 336200
rect 357600 330800 359300 336200
rect 359800 330800 360700 336200
rect 360800 330800 361100 336200
rect 361400 330800 363000 336200
rect 363500 330800 364500 336200
rect 364600 330800 364900 336200
rect 365200 330800 366800 336200
rect 367300 330800 368200 336200
rect 368300 330800 368600 336200
rect 368900 330800 370600 336200
rect 371100 330800 372000 336200
rect 372100 330800 372400 336200
rect 372700 330800 374300 336200
rect 374800 330800 375800 336200
rect 375900 330800 376200 336200
rect 376500 330800 378100 336200
rect 378600 330800 379500 336200
rect 379600 330800 379900 336200
rect 380200 330800 381800 336200
rect 382300 330800 383300 336200
rect 383400 330800 383700 336200
rect 384000 330800 385600 336200
rect 386100 330800 387100 336200
rect 387200 330800 387500 336200
rect 387800 330800 389400 336200
rect 389900 330800 390800 336200
rect 391000 330800 392200 336200
rect 392500 330800 394300 336200
rect 395800 330800 396800 336200
rect 397800 330800 400600 336200
rect 401800 330800 404900 336200
rect 405400 330800 406500 336200
rect 406600 330800 406900 336200
rect 407300 330800 408800 336200
rect 409300 330800 410300 336200
rect 410400 330800 410700 336200
rect 411000 330800 412600 336200
rect 413100 330800 414000 336200
rect 414100 330800 414400 336200
rect 414700 330800 416400 336200
rect 416900 330800 417800 336200
rect 417900 330800 418200 336200
rect 418500 330800 420100 336200
rect 420600 330800 421600 336200
rect 421700 330800 422000 336200
rect 422300 330800 423900 336200
rect 424400 330800 425300 336200
rect 425400 330800 425700 336200
rect 426000 330800 427600 336200
rect 428100 330800 429100 336200
rect 429200 330800 429500 336200
rect 429800 330800 431400 336200
rect 431900 330800 432800 336200
rect 432900 330800 433300 336200
rect 433600 330800 435200 336200
rect 435700 330800 436600 336200
rect 436700 330800 437000 336200
rect 437300 330800 438900 336200
rect 439400 330800 440400 336200
rect 440500 330800 440800 336200
rect 441100 330800 442700 336200
rect 443200 330800 444100 336200
rect 444200 330800 444600 336200
rect 444900 330800 446500 336200
rect 452600 330800 454000 336200
rect 454500 330800 455400 336200
rect 455500 330800 455800 336200
rect 456200 330800 457800 336200
rect 458300 330800 459200 336200
rect 459300 330800 459600 336200
rect 459900 330800 461500 336200
rect 462000 330800 463000 336200
rect 463100 330800 463400 336200
rect 463700 330800 465300 336200
rect 465800 330800 466800 336200
rect 467600 330800 472387 336200
rect 316853 330742 447000 330800
rect 452600 330742 472387 330800
rect 477987 330742 478200 336342
rect 316853 321813 317988 330742
rect 319000 323142 319295 328742
rect 324895 328600 478351 328742
rect 324895 323200 328200 328600
rect 329000 323200 330200 328600
rect 330300 323200 331600 328600
rect 332600 323200 333700 328600
rect 334000 323200 335400 328600
rect 336400 323200 337500 328600
rect 337800 323200 339200 328600
rect 340200 323200 340600 328600
rect 345800 323200 346700 328600
rect 347700 323200 348800 328600
rect 349100 323200 350400 328600
rect 351400 323200 352600 328600
rect 352900 323200 354200 328600
rect 355200 323200 356300 328600
rect 356600 323200 358000 328600
rect 359000 323200 360100 328600
rect 360400 323200 361700 328600
rect 362700 323200 363900 328600
rect 364200 323200 365500 328600
rect 366500 323200 367600 328600
rect 367900 323200 369200 328600
rect 370200 323200 371400 328600
rect 371700 323200 373000 328600
rect 374000 323200 375100 328600
rect 375400 323200 376800 328600
rect 377800 323200 378900 328600
rect 379200 323200 380600 328600
rect 381600 323200 382700 328600
rect 383000 323200 384300 328600
rect 385300 323200 386400 328600
rect 386700 323200 388100 328600
rect 389100 323200 390200 328600
rect 390500 323200 391300 328600
rect 391700 323200 392800 328600
rect 393800 323200 396100 328600
rect 396400 323200 398200 328600
rect 400000 323200 402300 328600
rect 403300 323200 403600 328600
rect 404600 323200 405700 328600
rect 406200 323200 407500 328600
rect 408500 323200 409700 328600
rect 410000 323200 411300 328600
rect 412300 323200 413400 328600
rect 413700 323200 415100 328600
rect 416100 323200 417200 328600
rect 417500 323200 418800 328600
rect 419800 323200 420900 328600
rect 421200 323200 422600 328600
rect 423600 323200 424700 328600
rect 425000 323200 426400 328600
rect 427400 323200 428500 328600
rect 428800 323200 430100 328600
rect 431100 323200 432300 328600
rect 432600 323200 433900 328600
rect 434900 323200 436000 328600
rect 436300 323200 437600 328600
rect 438600 323200 439800 328600
rect 440100 323200 441400 328600
rect 442400 323200 443500 328600
rect 443800 323200 445200 328600
rect 446200 323200 447300 328600
rect 447600 323200 448900 328600
rect 449900 323200 451100 328600
rect 451400 323200 452700 328600
rect 453700 323200 454800 328600
rect 455100 323200 456500 328600
rect 457500 323200 458600 328600
rect 458900 323200 460200 328600
rect 461200 323200 462400 328600
rect 462700 323200 464000 328600
rect 465000 323200 466100 328600
rect 466400 323200 467900 328600
rect 468600 323200 478351 328600
rect 324895 323142 478351 323200
rect 316853 320678 326140 321813
rect 472958 321527 473098 323142
rect 477488 321511 477628 323142
rect 321310 319704 321450 320678
rect 325840 319685 325980 320678
rect 37548 315630 38808 315756
rect 37548 314874 37674 315630
rect 38682 314874 38808 315630
rect 37548 314622 38808 314874
rect 37548 314496 80136 314622
rect 37548 313740 52668 314496
rect 54054 313740 58590 314496
rect 59346 313740 63756 314496
rect 65016 313740 68670 314496
rect 69426 313740 74592 314496
rect 80010 313740 80136 314496
rect 37548 313614 80136 313740
rect 35028 313488 36036 313614
rect 35028 312984 35154 313488
rect 35910 312984 36036 313488
rect 35028 312858 36036 312984
rect 42714 312858 42840 313614
rect 43218 312858 43344 313614
rect 42714 312732 43344 312858
rect 34146 311094 72450 311220
rect 34146 310212 34398 311094
rect 37044 310842 44100 311094
rect 37044 310338 42840 310842
rect 43218 310338 44100 310842
rect 37044 310212 44100 310338
rect 44352 310842 64512 311094
rect 44352 310338 50022 310842
rect 50400 310338 64512 310842
rect 44352 310212 64512 310338
rect 65394 310212 72450 311094
rect 34146 310086 72450 310212
rect 36328 309582 87822 309708
rect 36328 309078 50652 309582
rect 51282 309078 59346 309582
rect 36328 308826 59346 309078
rect 61362 308826 82278 309582
rect 87570 308826 87822 309582
rect 36328 308700 87822 308826
rect 54498 286272 80164 286412
rect 54498 285642 54936 286272
rect 55818 285642 57960 286272
rect 60354 285642 74592 286272
rect 80010 285642 80164 286272
rect 54498 285530 80164 285642
rect 48754 284886 87696 285012
rect 48754 284256 49266 284886
rect 50148 284256 82278 284886
rect 87570 284256 87696 284886
rect 48754 284130 87696 284256
rect 58401 247968 87822 248094
rect 58401 247086 58590 247968
rect 59220 247086 82278 247968
rect 87570 247086 87822 247968
rect 58401 246960 87822 247086
rect 60102 246330 60982 246456
rect 60102 245448 60228 246330
rect 60858 245448 60982 246330
rect 60102 243306 60982 245448
rect 63756 244692 87696 244818
rect 63756 243936 63882 244692
rect 64638 243936 82278 244692
rect 87570 243936 87696 244692
rect 63756 243810 87696 243936
rect 34272 243288 68670 243306
rect 34272 243180 44334 243288
rect 34272 242298 34398 243180
rect 37170 242298 44334 243180
rect 34272 242190 44334 242298
rect 44526 243180 68670 243288
rect 44526 242298 67284 243180
rect 67914 242298 68670 243180
rect 44526 242190 68670 242298
rect 34272 242172 68670 242190
rect 44636 241428 64372 242172
rect 65638 241794 67024 241920
rect 65638 241290 65764 241794
rect 66898 241290 67024 241794
rect 65638 241038 67024 241290
rect 65638 240912 80136 241038
rect 49644 239904 65268 240408
rect 65638 240156 74718 240912
rect 80010 240156 80136 240912
rect 65638 240030 80136 240156
rect 49644 239778 49770 239904
rect 51660 239778 65268 239904
rect 49644 239652 65268 239778
rect 64512 238896 65268 239652
rect 64512 238770 87696 238896
rect 64512 238014 82278 238770
rect 87570 238014 87696 238770
rect 64512 237888 87696 238014
rect 66276 233604 80136 233730
rect 66276 232596 66402 233604
rect 66654 232596 74718 233604
rect 80010 232596 80136 233604
rect 66276 232470 80136 232596
rect 72324 229320 87570 229446
rect 72324 228690 72450 229320
rect 73584 228690 82278 229320
rect 87444 228690 87570 229320
rect 72324 228564 87570 228690
rect 65268 226674 80010 226800
rect 65268 225792 65394 226674
rect 66528 225792 74718 226674
rect 79884 225792 80010 226674
rect 65268 225666 80010 225792
rect 72828 209538 87570 209664
rect 72828 208656 72954 209538
rect 73584 208656 82278 209538
rect 87444 208656 87570 209538
rect 72828 208530 87570 208656
rect 79254 207942 79758 208026
rect 79254 206980 79331 207942
rect 79685 206980 79758 207942
rect 79254 206892 79758 206980
rect 74306 205722 74654 205762
rect 74306 205038 74345 205722
rect 74614 205038 74654 205722
rect 74306 198976 74654 205038
rect 82278 200970 87696 201096
rect 82278 200340 82404 200970
rect 87570 200340 87696 200970
rect 82278 200214 87696 200340
rect 34272 198850 75096 198976
rect 34272 198094 34398 198850
rect 37170 198094 70812 198850
rect 71316 198094 75096 198850
rect 34272 197968 75096 198094
rect 49644 197316 87696 197442
rect 49644 197117 82278 197316
rect 49644 196869 49829 197117
rect 51830 196869 82278 197117
rect 49644 196812 82278 196869
rect 82152 196686 82278 196812
rect 87570 196686 87696 197316
rect 82152 196560 87696 196686
rect 68922 193032 87696 193158
rect 68922 192402 69048 193032
rect 69552 192402 82278 193032
rect 87570 192402 87696 193032
rect 68922 192276 87696 192402
rect 66024 190008 76482 190134
rect 66024 189252 66150 190008
rect 66780 189252 74592 190008
rect 76356 189252 76482 190008
rect 66024 189126 76482 189252
rect 65646 184212 80199 184338
rect 65646 183078 65772 184212
rect 66906 183078 74718 184212
rect 80010 183078 80199 184212
rect 65646 182952 80199 183078
rect 74844 167202 87696 167328
rect 74844 166446 74970 167202
rect 79632 166446 82278 167202
rect 87570 166446 87696 167202
rect 74844 166320 87696 166446
rect 79380 165312 80010 165438
rect 79380 164178 79506 165312
rect 79884 164178 80010 165312
rect 79380 164052 80010 164178
rect 70878 156752 71860 156878
rect 70878 156500 70964 156752
rect 71720 156500 71860 156752
rect 70878 155106 71860 156500
rect 71986 156792 87696 156870
rect 71986 156744 82278 156792
rect 71986 156492 72072 156744
rect 72828 156492 82278 156744
rect 87570 156492 87696 156792
rect 71986 156334 87696 156492
rect 71986 156333 72702 156334
rect 64638 155000 81648 155106
rect 34147 154980 81648 155000
rect 34147 154837 80892 154980
rect 34147 149710 34438 154837
rect 37165 154224 80892 154837
rect 81522 154224 81648 154980
rect 37165 154098 81648 154224
rect 37165 151956 66377 154098
rect 70812 153342 80136 153468
rect 70812 152964 70938 153342
rect 73710 152964 74718 153342
rect 80010 152964 80136 153342
rect 70812 152838 80136 152964
rect 37165 149710 59850 151956
rect 34147 149562 59850 149710
rect 60228 149562 66377 151956
rect 34147 149400 66377 149562
rect 60777 147250 66377 149400
rect 319090 147250 319230 151333
rect 321310 149844 321450 151300
rect 321000 149736 321600 149844
rect 321000 149336 321100 149736
rect 321500 149336 321600 149736
rect 321000 149236 321600 149336
rect 321000 148736 321600 148836
rect 321000 148336 321100 148736
rect 321500 148336 321600 148736
rect 321000 147250 321600 148336
rect 323620 147250 323760 151372
rect 60777 146412 98910 147250
rect 60777 142380 81270 146412
rect 81648 142380 98910 146412
rect 60777 141650 98910 142380
rect 99666 147212 118818 147250
rect 99666 141794 108864 147212
rect 114282 141794 118818 147212
rect 99666 141650 118818 141794
rect 119574 141650 138726 147250
rect 139482 141650 158634 147250
rect 159390 141650 178542 147250
rect 179298 141650 198450 147250
rect 199206 141650 218358 147250
rect 219114 141650 238266 147250
rect 239022 141650 258174 147250
rect 258930 141650 278082 147250
rect 278838 141650 297990 147250
rect 298746 147200 325000 147250
rect 298746 141800 319400 147200
rect 324800 141800 325000 147200
rect 298746 141650 325000 141800
rect 60777 139208 82144 139650
rect 60777 139198 69904 139208
rect 60777 135828 61910 139198
rect 60777 133560 60984 135828
rect 61362 134800 61910 135828
rect 65458 134800 69904 139198
rect 72582 134800 82144 139208
rect 61362 134050 82144 134800
rect 87744 139600 324173 139650
rect 87744 139340 311800 139600
rect 87744 139328 102056 139340
rect 87744 138432 89264 139328
rect 90720 138432 102056 139328
rect 87744 134800 102056 138432
rect 106736 134800 116382 139340
rect 87744 134658 116382 134800
rect 121206 139198 311800 139340
rect 121206 134658 209722 139198
rect 87744 134516 209722 134658
rect 214546 134516 311800 139198
rect 87744 134200 311800 134516
rect 317200 134200 324173 139600
rect 87744 134050 324173 134200
rect 61362 133560 66377 134050
rect 60777 131292 66377 133560
rect 60777 131040 62748 131292
rect 65646 131040 66377 131292
rect 60777 127008 66377 131040
rect 121464 131040 124956 131166
rect 74592 130662 80136 130788
rect 74592 130032 74718 130662
rect 80010 130032 80136 130662
rect 74592 129906 80136 130032
rect 121464 130032 121590 131040
rect 124866 130032 124956 131040
rect 121464 129906 124956 130032
rect 123956 128574 124956 129906
rect 125048 128574 126048 134050
rect 202734 132426 210974 133686
rect 202734 130032 202860 132426
rect 206010 130032 206136 132426
rect 209014 132174 210974 132426
rect 211170 132174 213130 134050
rect 275800 133700 276600 134050
rect 275800 133100 275900 133700
rect 276500 133100 276600 133700
rect 275800 133000 276600 133100
rect 275800 132300 276600 132400
rect 275800 131700 275900 132300
rect 276500 131700 276600 132300
rect 275800 131600 276600 131700
rect 276127 130664 276267 131600
rect 278347 130700 278487 134050
rect 282877 130700 283017 134050
rect 287407 130700 287547 134050
rect 291937 130700 292077 134050
rect 296467 130700 296607 134050
rect 300997 130700 301137 134050
rect 305527 130700 305667 134050
rect 310057 130700 310197 134050
rect 314587 130700 314727 134050
rect 319117 130700 319257 134050
rect 323647 130700 323787 134050
rect 60777 126630 61110 127008
rect 61866 126630 66377 127008
rect 34524 123000 35532 123102
rect 60777 123000 66377 126630
rect 34524 122976 50568 123000
rect 34524 117432 34650 122976
rect 35406 122460 50568 122976
rect 35406 117920 42618 122460
rect 47298 117920 50568 122460
rect 35406 117432 50568 117920
rect 34524 117400 50568 117432
rect 51352 122460 66377 123000
rect 51352 117920 61060 122460
rect 65740 117920 66377 122460
rect 51352 117400 66377 117920
rect 34524 116046 35532 117400
rect 34524 114912 34650 116046
rect 35406 114912 35532 116046
rect 34524 114786 35532 114912
rect 98784 111888 102816 112014
rect 74466 111636 80136 111762
rect 74466 110502 74592 111636
rect 80010 110502 80136 111636
rect 74466 110376 80136 110502
rect 98784 108612 98910 111888
rect 102690 108612 102816 111888
rect 98784 108486 102816 108612
rect 108738 110376 114282 110502
rect 108738 107100 108864 110376
rect 114156 107100 114282 110376
rect 108738 106974 114282 107100
rect 98784 84879 104328 85005
rect 98784 82782 98910 84879
rect 104202 82782 104328 84879
rect 98784 82656 104328 82782
rect 113148 75600 114030 75726
rect 40761 73332 103937 74113
rect 113148 73458 113274 75600
rect 113904 73458 114030 75600
rect 40761 73206 104328 73332
rect 40761 72586 98910 73206
rect 45469 71779 45609 72586
rect 49999 71779 50139 72586
rect 54529 71779 54669 72586
rect 59059 71779 59199 72586
rect 98784 71064 98910 72586
rect 96894 70938 98910 71064
rect 104202 71064 104328 73206
rect 113148 72072 114030 73458
rect 113148 71442 113274 72072
rect 113904 71442 114030 72072
rect 113148 71316 114030 71442
rect 123858 72828 140986 72954
rect 123858 71442 123984 72828
rect 128520 71442 136072 72828
rect 140860 71442 140986 72828
rect 123858 71316 140986 71442
rect 104202 70938 106344 71064
rect 96894 69426 97020 70938
rect 106218 69426 106344 70938
rect 96894 69300 106344 69426
rect 202734 58768 206136 130032
rect 475178 78607 475318 79670
rect 477488 79500 477628 79700
rect 477200 79400 477800 79500
rect 477200 79000 477300 79400
rect 477700 79000 477800 79400
rect 477200 78900 477800 79000
rect 479708 78607 479848 79660
rect 471132 78400 480110 78607
rect 471132 78000 477300 78400
rect 477700 78000 480110 78400
rect 471132 77028 480110 78000
rect 473724 75800 476475 77028
rect 472400 75600 478000 75800
rect 276127 64801 276267 65903
rect 280657 64801 280797 65903
rect 285187 64801 285327 65903
rect 289717 64801 289857 65903
rect 294247 64801 294387 65903
rect 298777 64801 298917 65903
rect 303307 64801 303447 65903
rect 307837 64801 307977 65903
rect 312367 64801 312507 65903
rect 316897 64801 317037 65903
rect 321427 64801 321567 65903
rect 274111 63290 324053 64801
rect 209014 58768 210974 62370
rect 211170 61614 213130 62370
rect 211170 59220 211302 61614
rect 213066 59220 213130 61614
rect 214194 61488 216154 62370
rect 274113 61488 283243 63290
rect 214194 61362 283248 61488
rect 214194 60228 268506 61362
rect 214200 59472 268506 60228
rect 283122 59472 283248 61362
rect 472400 61200 472600 75600
rect 477800 61200 478000 75600
rect 472400 61000 478000 61200
rect 214200 59346 283248 59472
rect 211170 59122 213130 59220
rect 285200 58768 300000 58800
rect 198934 58600 319295 58768
rect 34412 57800 40012 57920
rect 34400 57600 40012 57800
rect 34400 43200 34600 57600
rect 36200 43200 40012 57600
rect 198934 54266 285400 58600
rect 198934 53800 204646 54266
rect 198934 53168 199200 53800
rect 199000 51600 199200 53168
rect 204464 51600 204646 53800
rect 199000 51400 204646 51600
rect 205266 53800 285400 54266
rect 205266 51600 205440 53800
rect 210800 53400 285400 53800
rect 299800 53400 319295 58600
rect 210800 53168 319295 53400
rect 324895 53168 325200 58768
rect 210800 51600 211000 53168
rect 219134 52428 219275 53168
rect 223664 52428 223805 53168
rect 228194 52428 228335 53168
rect 232724 52428 232865 53168
rect 237254 52428 237395 53168
rect 241784 52428 241925 53168
rect 246314 52428 246455 53168
rect 250844 52428 250985 53168
rect 255374 52428 255515 53168
rect 259904 52428 260045 53168
rect 264434 52428 264575 53168
rect 268964 52428 269105 53168
rect 273494 52428 273635 53168
rect 278024 52428 278165 53168
rect 282554 52428 282695 53168
rect 287084 52428 287225 53168
rect 291614 52428 291755 53168
rect 296144 52428 296285 53168
rect 300674 52428 300815 53168
rect 305204 52428 305345 53168
rect 309734 52428 309875 53168
rect 314264 52428 314405 53168
rect 317800 52300 318600 53168
rect 317800 51700 317900 52300
rect 318500 51700 318600 52300
rect 317800 51600 318600 51700
rect 205266 51400 211000 51600
rect 316600 51100 318600 51200
rect 96138 50526 107604 50652
rect 96138 47754 96264 50526
rect 107478 47754 107604 50526
rect 316600 50500 317900 51100
rect 318500 50500 318600 51100
rect 316600 50400 318600 50500
rect 96138 47628 107604 47754
rect 34400 43000 40012 43200
rect 34412 40579 40012 43000
rect 59700 41785 60500 41800
rect 59192 41700 60500 41785
rect 43249 40579 43389 41563
rect 47779 40579 47919 41564
rect 52309 40579 52449 41556
rect 56839 40579 56979 41556
rect 59192 41540 59800 41700
rect 59700 41100 59800 41540
rect 60400 41100 60500 41700
rect 59700 41000 60500 41100
rect 59700 40579 60500 40600
rect 98784 40579 104384 47628
rect 321869 45793 323462 53168
rect 321869 45100 481596 45793
rect 321869 44500 480500 45100
rect 481100 44500 481596 45100
rect 321869 44200 481596 44500
rect 221354 42506 221494 43790
rect 225884 42506 226024 43790
rect 230414 42506 230554 43790
rect 234944 42515 235084 43790
rect 239474 42515 239614 43790
rect 244004 42515 244144 43790
rect 248534 42515 248674 43790
rect 253064 42515 253204 43790
rect 257594 42515 257734 43790
rect 262124 42515 262264 43790
rect 266654 42515 266794 43790
rect 271184 42515 271324 43790
rect 275714 42515 275854 43790
rect 280244 42515 280384 43790
rect 284774 42515 284914 43790
rect 289304 42515 289444 43790
rect 293834 42515 293974 43790
rect 298364 42515 298504 43790
rect 302894 42515 303034 43790
rect 307424 42515 307564 43790
rect 311954 42515 312094 43790
rect 316484 42519 316624 43790
rect 323794 43394 323934 44200
rect 328324 43394 328464 44200
rect 332854 43394 332994 44200
rect 337384 43394 337524 44200
rect 341914 43394 342054 44200
rect 346444 43394 346584 44200
rect 350974 43394 351114 44200
rect 355504 43394 355644 44200
rect 360034 43394 360174 44200
rect 364564 43394 364704 44200
rect 369094 43394 369234 44200
rect 373624 43394 373764 44200
rect 378154 43394 378294 44200
rect 382684 43394 382824 44200
rect 387214 43394 387354 44200
rect 391744 43394 391884 44200
rect 396274 43394 396414 44200
rect 400804 43394 400944 44200
rect 405334 43394 405474 44200
rect 409864 43394 410004 44200
rect 414394 43394 414534 44200
rect 418924 43394 419064 44200
rect 423454 43394 423594 44200
rect 427984 43394 428124 44200
rect 432514 43394 432654 44200
rect 437044 43394 437184 44200
rect 441574 43394 441714 44200
rect 446104 43394 446244 44200
rect 450634 43394 450774 44200
rect 455164 43394 455304 44200
rect 459694 43394 459834 44200
rect 464224 43394 464364 44200
rect 468754 43394 468894 44200
rect 473284 43394 473424 44200
rect 477814 43394 477954 44200
rect 480400 43700 481200 43800
rect 480400 43394 480500 43700
rect 480170 43100 480500 43394
rect 481100 43100 481200 43700
rect 480170 43033 481200 43100
rect 480400 43000 481200 43033
rect 315742 42515 317335 42519
rect 231600 42506 317388 42515
rect 218833 42400 317388 42506
rect 218833 42200 311800 42400
rect 218833 41154 231800 42200
rect 34412 40500 128772 40579
rect 34412 39900 59800 40500
rect 60400 40446 128772 40500
rect 60400 39900 123984 40446
rect 34412 35532 123984 39900
rect 128520 35532 128772 40446
rect 231600 37200 231800 41154
rect 246200 37200 311800 42200
rect 231600 37000 311800 37200
rect 317200 37000 317388 42400
rect 231600 36915 317388 37000
rect 34412 35400 128772 35532
rect 34412 34979 102400 35400
rect 102200 33800 102400 34979
rect 116800 34979 117298 35400
rect 116800 33800 117000 34979
rect 102200 33600 117000 33800
rect 315742 34238 317335 36915
rect 326014 34238 326154 34754
rect 330544 34238 330684 34754
rect 335074 34238 335214 34754
rect 339604 34238 339744 34754
rect 344134 34238 344274 34754
rect 348664 34238 348804 34754
rect 353194 34238 353334 34754
rect 357724 34238 357864 34754
rect 362254 34238 362394 34754
rect 366784 34238 366924 34754
rect 371314 34238 371454 34754
rect 375844 34238 375984 34754
rect 380374 34238 380514 34754
rect 384904 34238 385044 34754
rect 389434 34238 389574 34754
rect 393964 34238 394104 34754
rect 398494 34238 398634 34754
rect 403024 34238 403164 34754
rect 407554 34238 407694 34754
rect 412084 34238 412224 34754
rect 416614 34238 416754 34754
rect 421144 34238 421284 34754
rect 425674 34238 425814 34754
rect 430204 34238 430344 34754
rect 434734 34238 434874 34754
rect 439264 34238 439404 34754
rect 443794 34238 443934 34754
rect 448324 34238 448464 34754
rect 452854 34238 452994 34754
rect 457384 34238 457524 34754
rect 461914 34238 462054 34754
rect 466444 34238 466584 34754
rect 470974 34238 471114 34754
rect 475504 34238 475644 34754
rect 480034 34238 480174 34754
rect 315742 32645 480174 34238
<< viatpl >>
rect 319364 379520 324824 380634
rect 74544 366731 80144 372331
rect 82144 359131 87744 364731
rect 108864 359131 109620 364731
rect 128772 359131 129528 364731
rect 148680 359131 149436 364731
rect 168588 359131 169344 364731
rect 188496 359131 189252 364731
rect 208404 359131 209160 364731
rect 228312 359131 229068 364731
rect 248220 359131 248976 364731
rect 268128 359131 268884 364731
rect 288036 359131 288792 364731
rect 320796 365354 322407 365486
rect 322407 365354 322686 365486
rect 320796 364604 322686 365354
rect 447210 374222 452272 379208
rect 334600 360800 346000 362200
rect 35784 357588 37170 358470
rect 82278 335916 87570 336798
rect 472600 349200 477800 363600
rect 447000 336200 452600 336342
rect 447000 330800 447900 336200
rect 447900 330800 448000 336200
rect 448000 330800 448300 336200
rect 448300 330800 448600 336200
rect 448600 330800 450200 336200
rect 450200 330800 450700 336200
rect 450700 330800 451700 336200
rect 451700 330800 451800 336200
rect 451800 330800 452100 336200
rect 452100 330800 452400 336200
rect 452400 330800 452600 336200
rect 447000 330742 452600 330800
rect 472387 330742 477987 336342
rect 319295 323142 324895 328742
rect 340600 323200 341300 328600
rect 341300 323200 341600 328600
rect 341600 323200 342900 328600
rect 342900 323200 343900 328600
rect 343900 323200 345000 328600
rect 345000 323200 345300 328600
rect 345300 323200 345800 328600
rect 74592 313740 80010 314496
rect 35154 312984 35910 313488
rect 34398 310212 37044 311094
rect 82278 308826 87570 309582
rect 74592 285642 80010 286272
rect 82278 284256 87570 284886
rect 82278 247086 87570 247968
rect 82278 243936 87570 244692
rect 34398 242298 37170 243180
rect 74718 240156 80010 240912
rect 82278 238014 87570 238770
rect 74718 232596 80010 233604
rect 82278 228690 87444 229320
rect 74718 225792 79884 226674
rect 82278 208656 87444 209538
rect 79331 206980 79685 207942
rect 82404 200340 87570 200970
rect 34398 198094 37170 198850
rect 82278 196686 87570 197316
rect 82278 192402 87570 193032
rect 74592 189252 76356 190008
rect 74718 183078 80010 184212
rect 82278 166446 87570 167202
rect 79506 164178 79884 165312
rect 82278 156492 87570 156792
rect 34438 149710 37165 154837
rect 74718 152964 80010 153342
rect 98910 141650 99666 147250
rect 108864 141794 114282 147212
rect 118818 141650 119574 147250
rect 138726 141650 139482 147250
rect 158634 141650 159390 147250
rect 178542 141650 179298 147250
rect 198450 141650 199206 147250
rect 218358 141650 219114 147250
rect 238266 141650 239022 147250
rect 258174 141650 258930 147250
rect 278082 141650 278838 147250
rect 297990 141650 298746 147250
rect 319400 141800 324800 147200
rect 61910 134800 65458 139198
rect 69904 134800 72582 139208
rect 82144 134050 87744 139650
rect 102056 134800 106736 139340
rect 116382 134658 121206 139340
rect 209722 134516 214546 139198
rect 311800 134200 317200 139600
rect 74718 130032 80010 130662
rect 34650 117432 35406 122976
rect 42618 117920 47298 122460
rect 50568 117400 51352 123000
rect 61060 117920 65740 122460
rect 74592 110502 80010 111636
rect 98910 108612 102690 111888
rect 108864 107100 114156 110376
rect 98910 82782 104202 84879
rect 113274 73458 113904 75600
rect 98910 70938 104202 73206
rect 123984 71442 128520 72828
rect 98910 69552 104202 70938
rect 472600 61200 477800 75600
rect 319295 53168 324895 58768
rect 123984 35532 128520 40446
rect 311800 37000 317200 42400
<< metaltpl >>
rect 319295 380634 324895 380716
rect 319295 379520 319364 380634
rect 324824 379520 324895 380634
rect 74544 372331 80144 372600
rect 34243 358470 37262 358863
rect 34243 357588 35784 358470
rect 37170 357588 37262 358470
rect 34243 313488 37262 357588
rect 34243 312984 35154 313488
rect 35910 312984 37262 313488
rect 34243 311094 37262 312984
rect 34243 310212 34398 311094
rect 37044 310212 37262 311094
rect 34243 243180 37262 310212
rect 34243 242298 34398 243180
rect 37170 242298 37262 243180
rect 34243 198850 37262 242298
rect 34243 198094 34398 198850
rect 37170 198094 37262 198850
rect 34243 154837 37262 198094
rect 34243 149710 34438 154837
rect 37165 149710 37262 154837
rect 34243 149547 37262 149710
rect 74544 314496 80144 366731
rect 319295 365486 324895 379520
rect 447006 379208 452606 379484
rect 447006 375800 447210 379208
rect 74544 313740 74592 314496
rect 80010 313740 80144 314496
rect 74544 286272 80144 313740
rect 74544 285642 74592 286272
rect 80010 285642 80144 286272
rect 74544 241290 80144 285642
rect 82144 364731 87744 365000
rect 108864 364731 109620 364800
rect 87744 359778 108864 363750
rect 82144 336798 87744 359131
rect 128772 364731 129528 364800
rect 109620 359778 128772 363750
rect 108864 356600 109620 359131
rect 148680 364731 149436 364800
rect 129528 359778 148680 363750
rect 128772 356600 129528 359131
rect 168588 364731 169344 364800
rect 149436 359778 168588 363750
rect 148680 356600 149436 359131
rect 188496 364731 189252 364800
rect 169344 359778 188496 363750
rect 168588 356600 169344 359131
rect 208404 364731 209160 364800
rect 189252 359778 208404 363750
rect 188496 356600 189252 359131
rect 228312 364731 229068 364800
rect 209160 359778 228312 363750
rect 208404 356600 209160 359131
rect 248220 364731 248976 364800
rect 229068 359778 248220 363750
rect 228312 356600 229068 359131
rect 268128 364731 268884 364800
rect 248976 359778 268128 363750
rect 248220 356600 248976 359131
rect 288036 364731 288792 364800
rect 268884 359778 288036 363750
rect 268128 356600 268884 359131
rect 319295 364604 320796 365486
rect 322686 364604 324895 365486
rect 288792 359778 290294 363750
rect 288036 356600 288792 359131
rect 82144 335916 82278 336798
rect 87570 335916 87744 336798
rect 82144 309582 87744 335916
rect 82144 308826 82278 309582
rect 87570 308826 87744 309582
rect 82144 284886 87744 308826
rect 82144 284256 82278 284886
rect 87570 284256 87744 284886
rect 82144 247968 87744 284256
rect 82144 247086 82278 247968
rect 87570 247086 87744 247968
rect 82144 244692 87744 247086
rect 82144 243936 82278 244692
rect 87570 243936 87744 244692
rect 82144 241290 87744 243936
rect 74544 240912 80136 241290
rect 74544 240156 74718 240912
rect 80010 240156 80136 240912
rect 74544 239904 80136 240156
rect 82152 239904 87744 241290
rect 74544 233604 80144 239904
rect 74544 232596 74718 233604
rect 80010 232596 80144 233604
rect 74544 226674 80144 232596
rect 74544 225792 74718 226674
rect 79884 225792 80144 226674
rect 74544 207942 80144 225792
rect 74544 206980 79331 207942
rect 79685 206980 80144 207942
rect 74544 190008 80144 206980
rect 74544 189252 74592 190008
rect 76356 189252 80144 190008
rect 74544 184212 80144 189252
rect 74544 183078 74718 184212
rect 80010 183078 80144 184212
rect 74544 165312 80144 183078
rect 74544 164178 79506 165312
rect 79884 164178 80144 165312
rect 74544 153342 80144 164178
rect 74544 152964 74718 153342
rect 80010 152964 80144 153342
rect 61744 134800 61910 138996
rect 65458 134942 69904 139056
rect 35406 118204 38648 122176
rect 40152 114408 40936 124688
rect 50568 123000 51352 124600
rect 42478 118062 42618 122316
rect 47298 118062 50568 122316
rect 61744 122460 65298 134800
rect 74544 130662 80144 152964
rect 74544 130032 74718 130662
rect 80010 130032 80144 130662
rect 51352 118062 61060 122316
rect 74544 114408 80144 130032
rect 40152 112596 80144 114408
rect 82144 238770 87744 239904
rect 82144 238014 82278 238770
rect 87570 238014 87744 238770
rect 82144 229320 87744 238014
rect 82144 228690 82278 229320
rect 87444 228690 87744 229320
rect 82144 209538 87744 228690
rect 82144 208656 82278 209538
rect 87444 208656 87744 209538
rect 82144 200970 87744 208656
rect 82144 200340 82404 200970
rect 87570 200340 87744 200970
rect 82144 197316 87744 200340
rect 82144 196686 82278 197316
rect 87570 196686 87744 197316
rect 82144 193032 87744 196686
rect 82144 192402 82278 193032
rect 87570 192402 87744 193032
rect 82144 167202 87744 192402
rect 82144 166446 82278 167202
rect 87570 166446 87744 167202
rect 82144 156792 87744 166446
rect 82144 156492 82278 156792
rect 87570 156492 87744 156792
rect 82144 139650 87744 156492
rect 319295 328742 324895 364604
rect 447000 374222 447210 375800
rect 452272 374222 452606 379208
rect 447000 374004 452606 374222
rect 334400 362200 346200 362400
rect 334400 360800 334600 362200
rect 346000 360800 346200 362200
rect 334400 360600 346200 360800
rect 98910 147250 99666 148800
rect 97374 142744 98910 146432
rect 108735 147212 114335 147639
rect 108735 146432 108864 147212
rect 99666 142744 108864 146432
rect 98910 141600 99666 141650
rect 108735 141794 108864 142744
rect 114282 146432 114335 147212
rect 118818 147250 119574 148800
rect 114282 142744 118818 146432
rect 114282 141794 114335 142744
rect 87744 135084 102056 138914
rect 82144 119585 87744 134050
rect 82144 113985 104356 119585
rect 74544 111762 80144 112596
rect 74466 111636 80144 111762
rect 74466 110502 74592 111636
rect 80010 110502 80144 111636
rect 74466 110376 80144 110502
rect 74544 110348 80144 110376
rect 98756 111888 104356 113985
rect 98756 108612 98910 111888
rect 102690 108612 104356 111888
rect 12768 104160 16240 107184
rect 98756 84879 104356 108612
rect 98756 82782 98910 84879
rect 104202 82782 104356 84879
rect 98756 73206 104356 82782
rect 108735 110376 114335 141794
rect 138726 147250 139482 148800
rect 119574 142744 138726 146432
rect 118818 141600 119574 141650
rect 158634 147250 159390 148800
rect 139482 142744 158634 146432
rect 138726 141600 139482 141650
rect 178542 147250 179298 148800
rect 159390 142744 178542 146432
rect 158634 141600 159390 141650
rect 198450 147250 199200 148800
rect 218358 147250 219114 148800
rect 179298 142744 198450 146432
rect 178542 141600 179298 141650
rect 199206 142744 218358 146432
rect 238266 147250 239022 148800
rect 219114 142744 238266 146432
rect 198450 141600 199200 141650
rect 218358 141600 219114 141650
rect 258174 147250 258930 148800
rect 239022 142744 258174 146432
rect 238266 141600 239022 141650
rect 278082 147250 278838 148800
rect 258930 142744 278082 146432
rect 258174 141600 258930 141650
rect 297990 147250 298746 148800
rect 278838 142744 297990 146432
rect 278082 141600 278838 141650
rect 319295 147200 324895 323142
rect 340400 328600 346000 360600
rect 447000 336342 452600 374004
rect 447000 330600 452600 330742
rect 472387 363600 477987 365000
rect 472387 349200 472600 363600
rect 477800 349200 477987 363600
rect 472387 336342 477987 349200
rect 340400 323200 340600 328600
rect 345800 323200 346000 328600
rect 340400 323000 346000 323200
rect 319295 146432 319400 147200
rect 298746 142744 319400 146432
rect 297990 141600 298746 141650
rect 319295 141800 319400 142744
rect 324800 141800 324895 147200
rect 311695 139600 317295 140200
rect 121206 135084 209722 138772
rect 311695 138772 311800 139600
rect 214546 135084 311800 138772
rect 108735 107100 108864 110376
rect 114156 107100 114335 110376
rect 108735 75600 114335 107100
rect 108735 73458 113274 75600
rect 113904 73458 114335 75600
rect 108735 73329 114335 73458
rect 311695 134200 311800 135084
rect 317200 134200 317295 139600
rect 98756 71064 98910 73206
rect 104202 71064 104356 73206
rect 123858 72828 128646 72954
rect 123858 71442 123984 72828
rect 128520 71442 128646 72828
rect 12320 65296 16464 68544
rect 123858 40446 128646 71442
rect 123858 35532 123984 40446
rect 128520 35532 128646 40446
rect 311695 42515 317295 134200
rect 319295 58768 324895 141800
rect 319295 52600 324895 53168
rect 472387 75600 477987 330742
rect 472387 61200 472600 75600
rect 477800 61200 477987 75600
rect 472387 42515 477987 61200
rect 311695 42400 477987 42515
rect 311695 37000 311800 42400
rect 317200 37000 477987 42400
rect 311695 36915 477987 37000
rect 311695 36400 317295 36915
rect 472387 36906 477987 36915
rect 123858 35154 128646 35532
use dn_acpq8b  dn_acpq8b_32
timestamp 1567007490
transform 1 0 87517 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_33
timestamp 1567007490
transform 1 0 89111 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_34
timestamp 1567007490
transform 1 0 97709 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_35
timestamp 1567007490
transform 1 0 99303 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_28
timestamp 1567007490
transform 1 0 104317 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_29
timestamp 1567007490
transform 1 0 105911 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_30
timestamp 1567007490
transform 1 0 114509 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_31
timestamp 1567007490
transform 1 0 116103 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_24
timestamp 1567007490
transform 1 0 121117 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_25
timestamp 1567007490
transform 1 0 122711 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_26
timestamp 1567007490
transform 1 0 131309 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_27
timestamp 1567007490
transform 1 0 132903 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_20
timestamp 1567007490
transform 1 0 137917 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_21
timestamp 1567007490
transform 1 0 139511 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_22
timestamp 1567007490
transform 1 0 148109 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_23
timestamp 1567007490
transform 1 0 149703 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_16
timestamp 1567007490
transform 1 0 194717 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_17
timestamp 1567007490
transform 1 0 196311 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_18
timestamp 1567007490
transform 1 0 204909 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_19
timestamp 1567007490
transform 1 0 206503 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_12
timestamp 1567007490
transform 1 0 211517 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_13
timestamp 1567007490
transform 1 0 213111 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_14
timestamp 1567007490
transform 1 0 221709 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_15
timestamp 1567007490
transform 1 0 223303 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_8
timestamp 1567007490
transform 1 0 238317 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_9
timestamp 1567007490
transform 1 0 239911 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_10
timestamp 1567007490
transform 1 0 248509 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_11
timestamp 1567007490
transform 1 0 250103 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_4
timestamp 1567007490
transform 1 0 255117 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_5
timestamp 1567007490
transform 1 0 256711 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_6
timestamp 1567007490
transform 1 0 265309 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_7
timestamp 1567007490
transform 1 0 266903 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_1
timestamp 1567007490
transform 1 0 271917 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_0
timestamp 1567007490
transform 1 0 273511 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_2
timestamp 1567007490
transform 1 0 282109 0 1 381035
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_3
timestamp 1567007490
transform 1 0 283703 0 1 381013
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_36
timestamp 1567007490
transform 1 0 37117 0 1 378635
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_37
timestamp 1567007490
transform 1 0 38711 0 1 378613
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_38
timestamp 1567007490
transform 1 0 47309 0 1 378635
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_39
timestamp 1567007490
transform 1 0 48903 0 1 378613
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_40
timestamp 1567007490
transform 1 0 53917 0 1 378635
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_41
timestamp 1567007490
transform 1 0 55511 0 1 378613
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_42
timestamp 1567007490
transform 1 0 64109 0 1 378635
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_43
timestamp 1567007490
transform 1 0 65703 0 1 378613
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_44
timestamp 1567007490
transform 1 0 70717 0 1 378635
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_45
timestamp 1567007490
transform 1 0 72311 0 1 378613
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_46
timestamp 1567007490
transform 1 0 76709 0 1 378635
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_47
timestamp 1567007490
transform 1 0 78303 0 1 378613
box -209 -209 209 209
use cmm5t_q3aq8b  cmm5t_q3aq8b_0
timestamp 1565723183
transform 1 0 206692 0 1 372544
box -124505 -6480 124505 6480
use dn3_7x8jps  dn3_7x8jps_1
timestamp 1566571856
transform 1 0 470514 0 1 373214
box -314 -314 314 314
use dn_0f0tea  dn_0f0tea_3
timestamp 1566571856
transform 1 0 328914 0 1 365114
box -314 -314 314 314
use BU_3VX2  overtemp_level /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 321216 0 1 362544
box 0 0 672 896
use LS_3VX2  temp_level ~/design/ip/LS_3VX2/8/maglef
timestamp 1526911224
transform 1 0 317382 0 -1 360584
box 1992 -1320 3956 -168
use LS_3VX2  rcosc_ena_level
timestamp 1526911224
transform -1 0 67196 0 1 360840
box 1992 -1320 3956 -168
use BU_3VX2  rcosc_out_level
timestamp 1529525674
transform 1 0 63616 0 1 358064
box 0 0 672 896
use BU_3VX2  por_level
timestamp 1529525674
transform 1 0 64288 0 1 358064
box 0 0 672 896
use antenna_gtg92w  antenna_gtg92w_2
timestamp 1525700399
transform 1 0 272592 0 1 357476
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_3
timestamp 1525700399
transform 1 0 272844 0 1 357476
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_4
timestamp 1525700399
transform 1 0 273096 0 1 357476
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_5
timestamp 1525700399
transform 1 0 273348 0 1 357476
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_6
timestamp 1525700399
transform 1 0 273600 0 1 357476
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_7
timestamp 1525700399
transform 1 0 273852 0 1 357476
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_8
timestamp 1525700399
transform 1 0 274104 0 1 357476
box 0 0 140 140
use dn_acpq8b  dn_acpq8b_51
timestamp 1567007490
transform 0 -1 32855 1 0 338087
box -209 -209 209 209
use arcoc01_3v3  rcosc /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869549
transform 1 0 35406 0 1 337330
box 0 0 22400 20000
use aporc02_3v3  por /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869493
transform -1 0 64728 0 1 337452
box 0 0 5080 20000
use antenna_gtg92w  antenna_gtg92w_18
timestamp 1525700399
transform 1 0 89918 0 1 356050
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_17
timestamp 1525700399
transform 1 0 89918 0 1 355806
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_16
timestamp 1525700399
transform 1 0 89918 0 1 355562
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_15
timestamp 1525700399
transform 1 0 89918 0 1 355318
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_14
timestamp 1525700399
transform 1 0 89918 0 1 355074
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_13
timestamp 1525700399
transform 1 0 89918 0 1 354830
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_12
timestamp 1525700399
transform 1 0 89918 0 1 354586
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_11
timestamp 1525700399
transform 1 0 89918 0 1 354342
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_10
timestamp 1525700399
transform 1 0 89918 0 1 354098
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_9
timestamp 1525700399
transform 1 0 89918 0 1 353854
box 0 0 140 140
use dn_acpq8b  dn_acpq8b_50
timestamp 1567007490
transform 0 -1 32833 1 0 336605
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_52
timestamp 1567007490
transform 0 -1 32855 1 0 327895
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_53
timestamp 1567007490
transform 0 -1 32833 1 0 326301
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_48
timestamp 1567007490
transform 0 -1 32855 1 0 321287
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_49
timestamp 1567007490
transform 0 -1 32833 1 0 319805
box -209 -209 209 209
use acmpc01_3v3  comparator /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869319
transform -1 0 41836 0 -1 335248
box 0 0 5800 20000
use acsoc01_3v3  comp_bias /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869363
transform 1 0 43722 0 -1 335370
box 0 0 13600 20000
use acsoc02_3v3  opamp_bias /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869399
transform -1 0 68268 0 -1 335248
box 0 0 9300 20000
use dn_acpq8b  dn_acpq8b_54
timestamp 1567007490
transform 0 -1 32855 1 0 311095
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_55
timestamp 1567007490
transform 0 -1 32833 1 0 309501
box -209 -209 209 209
use AMUX4_3V  comp_ninput_mux ~/design/ip/AMUX4_3V/11/maglef
timestamp 1527118791
transform -1 0 47980 0 1 310738
box 5982 -1710 11512 2880
use AMUX4_3V  comp_pinput_mux
timestamp 1527118791
transform -1 0 55031 0 1 310746
box 5982 -1710 11512 2880
use BU_3VX2  comp_out_level
timestamp 1529525674
transform 1 0 62608 0 -1 313376
box 0 0 672 896
use AMUX2_3V  analog_out_mux ~/design/ip/AMUX2_3V/10/maglef
timestamp 1527162843
transform -1 0 62798 0 -1 311820
box 5694 -560 8904 2552
use LS_3VX2  comp_ena_level
timestamp 1526911224
transform -1 0 66452 0 -1 310619
box 1992 -1320 3956 -168
use LS_3VX2  opamp_ena_level
timestamp 1526911224
transform -1 0 68244 0 -1 310619
box 1992 -1320 3956 -168
use LS_3VX2  opamp_bias_ena_level
timestamp 1526911224
transform -1 0 70036 0 -1 310619
box 1992 -1320 3956 -168
use dn_acpq8b  dn_acpq8b_62
timestamp 1567007490
transform 0 -1 32599 1 0 304493
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_63
timestamp 1567007490
transform 0 -1 32577 1 0 302899
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_60
timestamp 1567007490
transform 0 -1 32599 1 0 294181
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_61
timestamp 1567007490
transform 0 -1 32577 1 0 292587
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_58
timestamp 1567007490
transform 0 -1 32615 1 0 288633
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_59
timestamp 1567007490
transform 0 -1 32593 1 0 287839
box -209 -209 209 209
use aopac01_3v3  opamp /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869437
transform -1 0 67928 0 -1 307798
box 0 0 30800 20000
use dn_acpq8b  dn_acpq8b_56
timestamp 1567007490
transform 0 -1 33155 1 0 277495
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_57
timestamp 1567007490
transform 0 -1 33133 1 0 275901
box -209 -209 209 209
use adacc01_3v3  dac /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869421
transform 0 -1 61942 1 0 244396
box 0 0 39116 23418
use AMUX4_3V  adc0_input_mux
timestamp 1527118791
transform 0 -1 69578 -1 0 240184
box 5982 -1710 11512 2880
use aadcc01_3v3  adc0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869217
transform 0 -1 72399 1 0 200236
box 0 0 39116 32500
use AMUX4_3V  adc1_input_mux
timestamp 1527118791
transform 0 -1 69704 -1 0 197248
box 5982 -1710 11512 2880
use aadcc01_3v3  adc1
timestamp 1513869217
transform 0 -1 72400 1 0 157414
box 0 0 39116 32500
use LOGIC1_3V  LOGIC1_3V_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 52691 0 1 147736
box 0 -80 560 976
use LOGIC1_3V  LOGIC1_3V_1
timestamp 1529525674
transform -1 0 53251 0 1 147736
box 0 -80 560 976
use LOGIC1_3V  LOGIC1_3V_2
timestamp 1529525674
transform -1 0 53811 0 1 147736
box 0 -80 560 976
use LOGIC1_3V  LOGIC1_3V_3
timestamp 1529525674
transform -1 0 54371 0 1 147736
box 0 -80 560 976
use ravenna_soc  ravenna_soc_0
timestamp 1567109375
transform 1 0 91098 0 1 148962
box -406 -394 225064 208282
use atmpc01_3v3  temp /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869651
transform -1 0 338908 0 -1 360047
box 0 0 18680 20000
use cmm5t_tqfh9t  cmm5t_tqfh9t_0
timestamp 1565723183
transform 1 0 444527 0 1 357522
box -27110 -15120 27110 15120
use dn_acpq8b  dn_acpq8b_68
timestamp 1567007490
transform 0 -1 477589 1 0 332463
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_69
timestamp 1567007490
transform 0 -1 477605 1 0 331037
box -209 -209 209 209
use cmm5t_g2pigg  cmm5t_g2pigg_0
timestamp 1565723183
transform 1 0 321520 0 1 235504
box -4460 -84240 4460 84240
use dn_0f0tea  dn_0f0tea_0
timestamp 1566571856
transform 1 0 321314 0 -1 148522
box -314 -314 314 314
use LOGIC0_3V  prog_ground_3 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 52030 0 -1 146999
box 0 0 560 896
use LOGIC0_3V  prog_ground_2
timestamp 1529525674
transform 1 0 52590 0 -1 146999
box 0 0 560 896
use LOGIC0_3V  prog_ground_1
timestamp 1529525674
transform 1 0 53150 0 -1 146999
box 0 0 560 896
use LOGIC0_3V  prog_ground_0
timestamp 1529525674
transform 1 0 53710 0 -1 146999
box 0 0 560 896
use ravenna_spi  ravenna_spi_0
timestamp 1567005482
transform 1 0 34160 0 1 124880
box -252 -336 24108 20972
use BU_3VX2  SCK_core_level
timestamp 1529525674
transform 1 0 61208 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_prod_id_level_7
timestamp 1529525674
transform 1 0 61880 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_prod_id_level_6
timestamp 1529525674
transform 1 0 62552 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_prod_id_level_5
timestamp 1529525674
transform 1 0 63224 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_prod_id_level_4
timestamp 1529525674
transform 1 0 63896 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_prod_id_level_3
timestamp 1529525674
transform 1 0 64568 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_prod_id_level_2
timestamp 1529525674
transform 1 0 65240 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_prod_id_level_1
timestamp 1529525674
transform 1 0 65912 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_prod_id_level_0
timestamp 1529525674
transform 1 0 66584 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_0
timestamp 1529525674
transform 1 0 67256 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_1
timestamp 1529525674
transform 1 0 67928 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_2
timestamp 1529525674
transform 1 0 68600 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_3
timestamp 1529525674
transform 1 0 69272 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_4
timestamp 1529525674
transform 1 0 69944 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_5
timestamp 1529525674
transform 1 0 70616 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_6
timestamp 1529525674
transform 1 0 71288 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_7
timestamp 1529525674
transform 1 0 71960 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_8
timestamp 1529525674
transform 1 0 72632 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_9
timestamp 1529525674
transform 1 0 73304 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_10
timestamp 1529525674
transform 1 0 73976 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mfgr_id_level_11
timestamp 1529525674
transform 1 0 74648 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mask_rev_level_0
timestamp 1529525674
transform 1 0 75320 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mask_rev_level_1
timestamp 1529525674
transform 1 0 75992 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mask_rev_level_2
timestamp 1529525674
transform 1 0 76664 0 -1 145320
box 0 0 672 896
use BU_3VX2  spi_mask_rev_level_3
timestamp 1529525674
transform 1 0 77336 0 -1 145320
box 0 0 672 896
use BU_3VX2  pass_thru_sck_level
timestamp 1529525674
transform 1 0 78008 0 -1 145320
box 0 0 672 896
use BU_3VX2  pass_thru_csb_level
timestamp 1529525674
transform 1 0 78680 0 -1 145320
box 0 0 672 896
use BU_3VX2  pass_thru_sdi_level
timestamp 1529525674
transform 1 0 79352 0 -1 145320
box 0 0 672 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 84394 0 -1 145656
box 0 -80 224 976
use IN_3VX2  IN_3VX2_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 84618 0 -1 145656
box 0 -80 448 976
use IN_3VX2  IN_3VX2_1
timestamp 1529525674
transform 1 0 85066 0 -1 145656
box 0 -80 448 976
use BU_3VX2  reg_ena_buf0
timestamp 1529525674
transform 1 0 85514 0 -1 145656
box 0 0 672 896
use BU_3VX2  reg_ena_buf1
timestamp 1529525674
transform 1 0 86186 0 -1 145656
box 0 0 672 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0
timestamp 1529525674
transform 1 0 86858 0 -1 145656
box 0 -80 224 976
use BU_3VX2  spi_config_level_7
timestamp 1529525674
transform 1 0 61768 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_config_level_6
timestamp 1529525674
transform 1 0 62440 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_config_level_5
timestamp 1529525674
transform 1 0 63112 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_config_level_4
timestamp 1529525674
transform 1 0 63784 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_config_level_3
timestamp 1529525674
transform 1 0 64456 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_config_level_2
timestamp 1529525674
transform 1 0 65128 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_config_level_1
timestamp 1529525674
transform 1 0 65800 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_config_level_0
timestamp 1529525674
transform 1 0 66472 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_irq_level
timestamp 1529525674
transform 1 0 67144 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_reg_enb_level
timestamp 1529525674
transform 1 0 67816 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_reg_ena_level
timestamp 1529525674
transform -1 0 69160 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_reset_level
timestamp 1529525674
transform 1 0 69160 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_pll_bypass_level
timestamp 1529525674
transform 1 0 69832 0 -1 135800
box 0 0 672 896
use BU_3VX2  pll_vco_ena_level
timestamp 1529525674
transform 1 0 70504 0 -1 135800
box 0 0 672 896
use BU_3VX2  pll_cp_ena_level
timestamp 1529525674
transform 1 0 71176 0 -1 135800
box 0 0 672 896
use BU_3VX2  pll_bias_ena_level
timestamp 1529525674
transform 1 0 71848 0 -1 135800
box 0 0 672 896
use BU_3VX2  spi_xtal_ena_level
timestamp 1529525674
transform 1 0 72520 0 -1 135800
box 0 0 672 896
use BU_3VX2  pll_vco_in_level
timestamp 1529525674
transform 1 0 73192 0 -1 135800
box 0 0 672 896
use BU_3VX2  pll_trim_level_3
timestamp 1529525674
transform 1 0 73864 0 -1 135800
box 0 0 672 896
use BU_3VX2  pll_trim_level_2
timestamp 1529525674
transform 1 0 74536 0 -1 135800
box 0 0 672 896
use BU_3VX2  pll_trim_level_1
timestamp 1529525674
transform 1 0 75208 0 -1 135800
box 0 0 672 896
use BU_3VX2  pll_trim_level_0
timestamp 1529525674
transform 1 0 75880 0 -1 135800
box 0 0 672 896
use BU_3VX2  pass_thru_level
timestamp 1529525674
transform 1 0 76552 0 -1 135800
box 0 0 672 896
use BU_3VX2  tm_nvcp_level_0
timestamp 1529525674
transform 1 0 77224 0 -1 135800
box 0 0 672 896
use BU_3VX2  tm_nvcp_level_1
timestamp 1529525674
transform 1 0 77896 0 -1 135800
box 0 0 672 896
use BU_3VX2  tm_nvcp_level_2
timestamp 1529525674
transform 1 0 78568 0 -1 135800
box 0 0 672 896
use BU_3VX2  tm_nvcp_level_3
timestamp 1529525674
transform 1 0 79240 0 -1 135800
box 0 0 672 896
use LOGIC0_3V  spi_config_zero_7
timestamp 1529525674
transform 1 0 61662 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  spi_config_zero_6
timestamp 1529525674
transform 1 0 62222 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  spi_config_zero_5
timestamp 1529525674
transform 1 0 62782 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  spi_config_zero_4
timestamp 1529525674
transform 1 0 63342 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  spi_config_zero_3
timestamp 1529525674
transform 1 0 63902 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  spi_config_zero_2
timestamp 1529525674
transform 1 0 64462 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  spi_config_zero_1
timestamp 1529525674
transform 1 0 65022 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  spi_config_zero_0
timestamp 1529525674
transform 1 0 65582 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  ground_digital
timestamp 1529525674
transform 1 0 66142 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_0
timestamp 1529525674
transform 1 0 66702 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_1
timestamp 1529525674
transform 1 0 67262 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_2
timestamp 1529525674
transform 1 0 67822 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_3
timestamp 1529525674
transform 1 0 68382 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_4
timestamp 1529525674
transform 1 0 68942 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_5
timestamp 1529525674
transform 1 0 69502 0 -1 133560
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_6
timestamp 1529525674
transform 1 0 70062 0 -1 133560
box 0 0 560 896
use LS_3VX2  pass_thru_sdo_level
timestamp 1526911224
transform -1 0 62274 0 -1 130015
box 1992 -1320 3956 -168
use LS_3VX2  spi_trap_level
timestamp 1526911224
transform -1 0 64066 0 -1 130015
box 1992 -1320 3956 -168
use LOGIC1  vdd_digital /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS
timestamp 1529525608
transform 1 0 58967 0 1 126596
box 0 0 252 976
use DFRX2  clock_div2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS
timestamp 1529525608
transform 1 0 62838 0 1 110948
box 0 -80 2520 1056
use DFRX2  clock_div4
timestamp 1529525608
transform 1 0 65358 0 1 110948
box 0 -80 2520 1056
use DFRX2  clock_div8
timestamp 1529525608
transform 1 0 67878 0 1 110948
box 0 -80 2520 1056
use BU_3VX2  xtal_out_level
timestamp 1529525674
transform 1 0 61440 0 1 108151
box 0 0 672 896
use BUX4  BUX4_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS
timestamp 1529525608
transform 1 0 63356 0 1 108168
box 0 -80 1008 1056
use BUX4  BUX4_0
timestamp 1529525608
transform 1 0 68122 0 1 108168
box 0 -80 1008 1056
use BUX12  BUX12_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS
timestamp 1529525608
transform 1 0 69130 0 1 108168
box 0 -80 2520 1056
use AMUX2_3V  vco_in_mux
timestamp 1527162843
transform -1 0 95592 0 -1 109960
box 5694 -560 8904 2552
use apllc03_1v8  pll /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_1V8
timestamp 1513868860
transform 1 0 38432 0 1 74948
box 0 0 54156 31048
use acsoc04_1v8  pll_bias /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_1V8
timestamp 1513868641
transform -1 0 107911 0 1 84085
box 0 0 13200 22000
use XNVR_136X32P128_VD01  nvram ~/design/ip/XNVR_136X32P128_VD01/1/maglef
timestamp 1555448905
transform 1 0 119923 0 -1 128630
box 0 0 81772 52856
use antenna_gtg92w  antenna_gtg92w_1
timestamp 1525700399
transform 1 0 120144 0 1 72780
box 0 0 140 140
use antenna_gtg92w  antenna_gtg92w_0
timestamp 1525700399
transform 1 0 120142 0 1 72488
box 0 0 140 140
use cmm5t_plguac  cmm5t_plguac_0
timestamp 1565723183
transform 1 0 50209 0 1 56660
box -8990 -15120 8990 15120
use LS_3VX2  bg_ena_level
timestamp 1526911224
transform 1 0 113816 0 -1 70896
box 1992 -1320 3956 -168
use markings  markings_0 markings
timestamp 1555546719
transform 1 0 129298 0 1 -172033
box -69538 220921 -57665 242943
use abgpc01_3v3  bandgap /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1513869238
transform -1 0 130818 0 -1 70160
box 0 0 58208 20000
use XCPF_136X32DP128_VD03  nvram_cp ~/design/ip/XCPF_136X32DP128_VD03/1/maglef
timestamp 1555448811
transform 1 0 207842 0 -1 132181
box 0 0 64252 69857
use dn3_7x8jps  dn3_7x8jps_0
timestamp 1566571856
transform 1 0 276200 0 1 131956
box -314 -314 314 314
use cmm5t_jqtkwo  cmm5t_jqtkwo_0
timestamp 1565723183
transform 1 0 298942 0 1 98300
box -24845 -32400 24845 32400
use cmm5t_7yf5ef  cmm5t_7yf5ef_0
timestamp 1565723183
transform 1 0 266864 0 1 48108
box -49760 -4320 49760 4320
use dn_0f0tea  dn_0f0tea_1
timestamp 1566571856
transform 1 0 318214 0 1 52014
box -314 -314 314 314
use XSPRAMBLP_4096X32_M8P  XSPRAMBLP_4096X32_M8P_0 ~/design/ip/XSPRAMBLP_4096X32_M8P/1/maglef
timestamp 1562789036
transform -1 0 468681 0 -1 316496
box -120 0 140671 269755
use dn_acpq8b  dn_acpq8b_70
timestamp 1567007490
transform 0 -1 477589 1 0 315663
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_71
timestamp 1567007490
transform 0 -1 477605 1 0 314237
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_72
timestamp 1567007490
transform 0 -1 477589 1 0 298863
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_73
timestamp 1567007490
transform 0 -1 477605 1 0 297437
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_74
timestamp 1567007490
transform 0 -1 477589 1 0 225263
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_75
timestamp 1567007490
transform 0 -1 477605 1 0 223837
box -209 -209 209 209
use cmm5t_8etd0t  cmm5t_8etd0t_0
timestamp 1565723183
transform 1 0 475388 0 1 200580
box -4460 -120960 4460 120960
use dn_acpq8b  dn_acpq8b_66
timestamp 1567007490
transform 0 -1 481417 1 0 134997
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_67
timestamp 1567007490
transform 0 -1 481433 1 0 133571
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_64
timestamp 1567007490
transform 0 -1 481417 1 0 118197
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_65
timestamp 1567007490
transform 0 -1 481433 1 0 116771
box -209 -209 209 209
use dn_0f0tea  dn_0f0tea_2
timestamp 1566571856
transform 1 0 477514 0 1 79214
box -314 -314 314 314
use dn_0f0tea  dn_0f0tea_4
timestamp 1566571856
transform 1 0 480814 0 1 44814
box -314 -314 314 314
use dn3_7x8jps  dn3_7x8jps_2
timestamp 1566571856
transform 1 0 60114 0 1 40214
box -314 -314 314 314
use cmm5t_yvxjnn  cmm5t_yvxjnn_0
timestamp 1565723183
transform 1 0 400969 0 1 39074
box -79205 -4320 79205 4320
use dn_acpq8b  dn_acpq8b_86
timestamp 1567007490
transform 1 0 310947 0 -1 32821
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_87
timestamp 1567007490
transform 1 0 312373 0 -1 32805
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_84
timestamp 1567007490
transform 1 0 327747 0 -1 32821
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_85
timestamp 1567007490
transform 1 0 329173 0 -1 32805
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_82
timestamp 1567007490
transform 1 0 364547 0 -1 32821
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_83
timestamp 1567007490
transform 1 0 365973 0 -1 32805
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_80
timestamp 1567007490
transform 1 0 381347 0 -1 32821
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_81
timestamp 1567007490
transform 1 0 382773 0 -1 32805
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_78
timestamp 1567007490
transform 1 0 398147 0 -1 32821
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_79
timestamp 1567007490
transform 1 0 399573 0 -1 32805
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_77
timestamp 1567007490
transform 1 0 414947 0 -1 32821
box -209 -209 209 209
use dn_acpq8b  dn_acpq8b_76
timestamp 1567007490
transform 1 0 416373 0 -1 32805
box -209 -209 209 209
use ravenna_padframe  ravenna_padframe_0
timestamp 1567010579
transform 1 0 126673 0 1 79633
box -126673 -79633 387927 333967
<< labels >>
flabel metal2 60032 148848 60032 148848 0 FreeSans 640 90 0 0 pass_thru_sdo_lv
flabel metal2 61824 148848 61824 148848 0 FreeSans 640 90 0 0 trap_lv
flabel metal2 77056 148848 77056 148848 0 FreeSans 640 90 0 0 pass_thru_reset_lv
flabel metal2 76384 148848 76384 148848 0 FreeSans 640 90 0 0 pll_trim_0_lv
flabel metal2 75712 148848 75712 148848 0 FreeSans 640 90 0 0 pll_trim_1_lv
flabel metal2 75040 148848 75040 148848 0 FreeSans 640 90 0 0 pll_trim_2_lv
flabel metal2 74368 148848 74368 148848 0 FreeSans 640 90 0 0 pll_trim_3_lv
flabel metal2 73696 148848 73696 148848 0 FreeSans 640 90 0 0 pll_vco_in_lv
flabel metal2 73024 148848 73024 148848 0 FreeSans 640 90 0 0 spi_xtal_ena_lv
flabel metal2 72352 148848 72352 148848 0 FreeSans 640 90 0 0 pll_bias_ena_lv
flabel metal2 71680 148848 71680 148848 0 FreeSans 640 90 0 0 pll_cp_ena_lv
flabel metal2 71008 148848 71008 148848 0 FreeSans 640 90 0 0 pll_vco_ena_lv
flabel metal2 70336 148848 70336 148848 0 FreeSans 640 90 0 0 pll_bypass_lv
flabel metal2 69664 148848 69664 148848 0 FreeSans 640 90 0 0 spi_reset_lv
flabel metal2 68880 148848 68880 148848 0 FreeSans 640 90 0 0 spi_reg_ena_lv
flabel metal2 67872 148848 67872 148848 0 FreeSans 640 90 0 0 spi_irq_lv
flabel metal2 67200 148848 67200 148848 0 FreeSans 640 90 0 0 config_0_lv
flabel metal2 66528 148848 66528 148848 0 FreeSans 640 90 0 0 config_1_lv
flabel metal2 65856 148848 65856 148848 0 FreeSans 640 90 0 0 config_2_lv
flabel metal2 65184 148848 65184 148848 0 FreeSans 640 90 0 0 config_3_lv
flabel metal2 64512 148848 64512 148848 0 FreeSans 640 90 0 0 config_4_lv
flabel metal2 63840 148848 63840 148848 0 FreeSans 640 90 0 0 config_5_lv
flabel metal2 63168 148848 63168 148848 0 FreeSans 640 90 0 0 config_6_lv
flabel metal2 62496 148848 62496 148848 0 FreeSans 640 90 0 0 config_7_lv
flabel metal2 79184 148848 79184 148848 0 FreeSans 640 90 0 0 pass_thru_csb_lv
flabel metal2 78512 148848 78512 148848 0 FreeSans 640 90 0 0 pass_thru_sck_lv
flabel metal2 79856 148848 79856 148848 0 FreeSans 640 90 0 0 pass_thru_sdi_lv
flabel metal2 77840 148848 77840 148848 0 FreeSans 640 90 0 0 mask_rev_3_lv
flabel metal2 77168 148848 77168 148848 0 FreeSans 640 90 0 0 mask_rev_2_lv
flabel metal2 76496 148848 76496 148848 0 FreeSans 640 90 0 0 mask_rev_1_lv
flabel metal2 75824 148848 75824 148848 0 FreeSans 640 90 0 0 mask_rev_0_lv
flabel metal2 75152 148848 75152 148848 0 FreeSans 640 90 0 0 mfgr_id_11_lv
flabel metal2 74480 148848 74480 148848 0 FreeSans 640 90 0 0 mfgr_id_10_lv
flabel metal2 73808 148848 73808 148848 0 FreeSans 640 90 0 0 mfgr_id_9_lv
flabel metal2 73136 148848 73136 148848 0 FreeSans 640 90 0 0 mfgr_id_8_lv
flabel metal2 72464 148848 72464 148848 0 FreeSans 640 90 0 0 mfgr_id_7_lv
flabel metal2 71792 148848 71792 148848 0 FreeSans 640 90 0 0 mfgr_id_6_lv
flabel metal2 71120 148848 71120 148848 0 FreeSans 640 90 0 0 mfgr_id_5_lv
flabel metal2 70448 148848 70448 148848 0 FreeSans 640 90 0 0 mfgr_id_4_lv
flabel metal2 69776 148848 69776 148848 0 FreeSans 640 90 0 0 mfgr_id_3_lv
flabel metal2 69104 148848 69104 148848 0 FreeSans 640 90 0 0 mfgr_id_2_lv
flabel metal2 68432 148848 68432 148848 0 FreeSans 640 90 0 0 mfgr_id_1_lv
flabel metal2 67760 148848 67760 148848 0 FreeSans 640 90 0 0 mfgr_id_0_lv
flabel metal2 67088 148848 67088 148848 0 FreeSans 640 90 0 0 prod_id_0_lv
flabel metal2 66416 148848 66416 148848 0 FreeSans 640 90 0 0 prod_id_1_lv
flabel metal2 65744 148848 65744 148848 0 FreeSans 640 90 0 0 prod_id_2_lv
flabel metal2 65072 148848 65072 148848 0 FreeSans 640 90 0 0 prod_id_3_lv
flabel metal2 64400 148848 64400 148848 0 FreeSans 640 90 0 0 prod_id_4_lv
flabel metal2 63728 148848 63728 148848 0 FreeSans 640 90 0 0 prod_id_5_lv
flabel metal2 63056 148848 63056 148848 0 FreeSans 640 90 0 0 prod_id_6_lv
flabel metal2 62384 148848 62384 148848 0 FreeSans 640 90 0 0 prod_id_7_lv
flabel metal2 396144 336354 396144 336354 0 FreeSans 1008 90 0 0 cen
rlabel metal2 52500 123620 52556 123676 8 pll_trim[0]
rlabel metal2 56868 146692 56924 146748 6 mask_rev_in[3]
rlabel metal2 56644 146692 56700 146748 6 mask_rev_in[2]
rlabel metal2 55524 146692 55580 146748 6 mask_rev_in[1]
rlabel metal2 47236 146132 47292 146188 6 mask_rev_in[0]
rlabel metal2 44324 123620 44380 123676 8 pass_thru_reset
rlabel metal2 48916 123620 48972 123676 8 tm_nvcp[3]
rlabel metal2 51828 123620 51884 123676 8 tm_nvcp[2]
rlabel metal2 52052 123620 52108 123676 8 tm_nvcp[1]
rlabel metal2 52276 123620 52332 123676 8 tm_nvcp[0]
rlabel metal2 56308 123620 56364 123676 8 pll_trim[3]
rlabel metal2 53284 123620 53340 123676 8 pll_trim[2]
rlabel metal2 52724 123620 52780 123676 8 pll_trim[1]
flabel metal2 315098 359628 315154 359684 6 FreeSans 480 90 0 0 spi_master_sdoenb
flabel metal2 315854 359628 315910 359684 6 FreeSans 480 90 0 0 spi_master_sdo
flabel metal2 314846 359628 314902 359684 6 FreeSans 480 90 0 0 spi_master_sdi
flabel metal2 315350 359628 315406 359684 6 FreeSans 480 90 0 0 spi_master_sck
flabel metal2 315602 359628 315658 359684 6 FreeSans 480 90 0 0 spi_master_csb
flabel metal2 309554 359628 309610 359684 6 FreeSans 480 90 0 0 sda_padoeb
flabel metal2 309806 359628 309862 359684 6 FreeSans 480 90 0 0 sda_pad_o
flabel metal2 310058 359628 310114 359684 6 FreeSans 480 90 0 0 sda_pad_i
flabel metal2 309302 359628 309358 359684 6 FreeSans 480 90 0 0 scl_padoeb
flabel metal2 314090 359628 314146 359684 6 FreeSans 480 90 0 0 gpio_in[0]
flabel metal2 313838 359628 313894 359684 6 FreeSans 480 90 0 0 gpio_in[1]
flabel metal2 313586 359628 313642 359684 6 FreeSans 480 90 0 0 gpio_in[2]
flabel metal2 313334 359628 313390 359684 6 FreeSans 480 90 0 0 gpio_in[3]
flabel metal2 313082 359628 313138 359684 6 FreeSans 480 90 0 0 gpio_in[4]
flabel metal2 312830 359628 312886 359684 6 FreeSans 480 90 0 0 gpio_in[5]
flabel metal2 312578 359628 312634 359684 6 FreeSans 480 90 0 0 gpio_in[6]
flabel metal2 312326 359628 312382 359684 6 FreeSans 480 90 0 0 gpio_in[7]
flabel metal2 312074 359628 312130 359684 6 FreeSans 480 90 0 0 gpio_in[8]
flabel metal2 311822 359628 311878 359684 6 FreeSans 480 90 0 0 gpio_in[9]
flabel metal2 311570 359628 311626 359684 6 FreeSans 480 90 0 0 gpio_in[10]
flabel metal2 311318 359628 311374 359684 6 FreeSans 480 90 0 0 gpio_in[11]
flabel metal2 311066 359628 311122 359684 6 FreeSans 480 90 0 0 gpio_in[12]
flabel metal2 310814 359628 310870 359684 6 FreeSans 480 90 0 0 gpio_in[13]
flabel metal2 310562 359628 310618 359684 6 FreeSans 480 90 0 0 gpio_in[14]
flabel metal2 310310 359628 310366 359684 6 FreeSans 480 90 0 0 gpio_in[15]
flabel metal2 292040 359628 292096 359684 6 FreeSans 480 90 0 0 scl_pad_i
flabel metal2 292292 359628 292348 359684 6 FreeSans 480 90 0 0 scl_pad_o
flabel metal2 273644 359628 273700 359684 6 FreeSans 480 90 0 0 adc0_clk
flabel metal2 273896 359628 273952 359684 6 FreeSans 480 90 0 0 adc0_convert
flabel metal2 275408 359628 275464 359684 6 FreeSans 480 90 0 0 adc0_done
flabel metal2 274148 359628 274204 359684 6 FreeSans 480 90 0 0 adc0_ena
flabel metal2 272888 359628 272944 359684 6 FreeSans 480 90 0 0 adc1_clk
flabel metal2 273140 359628 273196 359684 6 FreeSans 480 90 0 0 adc1_convert
flabel metal2 275156 359628 275212 359684 6 FreeSans 480 90 0 0 adc1_done
flabel metal2 273392 359628 273448 359684 6 FreeSans 480 90 0 0 adc1_ena
flabel metal2 272384 359628 272440 359684 6 FreeSans 480 90 0 0 analog_out_sel
flabel metal2 271628 359628 271684 359684 6 FreeSans 480 90 0 0 bg_ena
flabel metal2 271376 359628 271432 359684 6 FreeSans 480 90 0 0 comp_ena
flabel metal2 274400 359628 274456 359684 6 FreeSans 480 90 0 0 comp_in
flabel metal2 272636 359628 272692 359684 6 FreeSans 480 90 0 0 dac_ena
flabel metal2 271880 359628 271936 359684 6 FreeSans 480 90 0 0 opamp_bias_ena
flabel metal2 272132 359628 272188 359684 6 FreeSans 480 90 0 0 opamp_ena
flabel metal2 274904 359628 274960 359684 6 FreeSans 480 90 0 0 overtemp
flabel metal2 270872 359628 270928 359684 6 FreeSans 480 90 0 0 overtemp_ena
flabel metal2 271124 359628 271180 359684 6 FreeSans 480 90 0 0 rcosc_ena
flabel metal2 274652 359628 274708 359684 6 FreeSans 480 90 0 0 rcosc_in
flabel metal2 270620 359628 270676 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[11]
flabel metal2 270368 359628 270424 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[10]
flabel metal2 270116 359628 270172 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[9]
flabel metal2 269864 359628 269920 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[8]
flabel metal2 269612 359628 269668 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[7]
flabel metal2 269360 359628 269416 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[6]
flabel metal2 269108 359628 269164 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[5]
flabel metal2 268856 359628 268912 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[4]
flabel metal2 268604 359628 268660 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[3]
flabel metal2 268352 359628 268408 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[2]
flabel metal2 266966 359628 267022 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[1]
flabel metal2 241514 359628 241570 359684 6 FreeSans 480 90 0 0 spi_ro_mfgr_id[0]
flabel metal2 230048 359628 230104 359684 6 FreeSans 480 90 0 0 spi_ro_pll_trim[1]
flabel metal2 229796 359628 229852 359684 6 FreeSans 480 90 0 0 spi_ro_pll_trim[2]
flabel metal2 232694 359628 232750 359684 6 FreeSans 480 90 0 0 spi_ro_pll_trim[0]
flabel metal2 232946 359628 233002 359684 6 FreeSans 480 90 0 0 comp_pinputsrc[0]
flabel metal2 233198 359628 233254 359684 6 FreeSans 480 90 0 0 comp_pinputsrc[1]
flabel metal2 199304 359628 199360 359684 6 FreeSans 480 90 0 0 comp_ninputsrc[1]
flabel metal2 206864 359628 206920 359684 6 FreeSans 480 90 0 0 comp_ninputsrc[0]
flabel metal2 209258 359628 209314 359684 6 FreeSans 480 90 0 0 spi_ro_pll_trim[3]
flabel metal2 202832 147348 202888 147404 8 FreeSans 480 90 0 0 xtal_in
flabel metal2 202580 147348 202636 147404 8 FreeSans 480 90 0 0 pll_clk
flabel metal2 203084 147348 203140 147404 8 FreeSans 480 90 0 0 flash_io3_do
flabel metal2 203336 147348 203392 147404 8 FreeSans 480 90 0 0 flash_io2_do
flabel metal2 203588 147348 203644 147404 8 FreeSans 480 90 0 0 flash_io1_do
flabel metal2 203840 147348 203896 147404 8 FreeSans 480 90 0 0 flash_io0_do
flabel metal2 201194 147348 201250 147404 8 FreeSans 480 90 0 0 ext_clk_sel
flabel metal2 202328 147348 202384 147404 8 FreeSans 480 90 0 0 ext_clk
flabel metal2 293930 146738 293986 146794 8 FreeSans 480 90 0 0 flash_clk_oeb
flabel metal2 293678 146738 293734 146794 8 FreeSans 480 90 0 0 flash_csb_oeb
flabel metal2 294434 146738 294490 146794 8 FreeSans 480 90 0 0 flash_io0_di
flabel metal2 293426 146738 293482 146794 8 FreeSans 480 90 0 0 flash_io0_oeb
flabel metal2 294686 146738 294742 146794 8 FreeSans 480 90 0 0 flash_io1_di
flabel metal2 293174 146738 293230 146794 8 FreeSans 480 90 0 0 flash_io1_oeb
flabel metal2 294938 146738 294994 146794 8 FreeSans 480 90 0 0 flash_io2_di
flabel metal2 295190 146738 295246 146794 8 FreeSans 480 90 0 0 flash_io3_di
flabel metal2 306026 146738 306082 146794 8 FreeSans 480 90 0 0 nvram_addr[7]
flabel metal2 306278 146738 306334 146794 8 FreeSans 480 90 0 0 nvram_addr[6]
flabel metal2 306530 146738 306586 146794 8 FreeSans 480 90 0 0 nvram_addr[5]
flabel metal2 306782 146738 306838 146794 8 FreeSans 480 90 0 0 nvram_addr[4]
flabel metal2 307034 146738 307090 146794 8 FreeSans 480 90 0 0 nvram_addr[3]
flabel metal2 307286 146738 307342 146794 8 FreeSans 480 90 0 0 nvram_addr[2]
flabel metal2 307538 146738 307594 146794 8 FreeSans 480 90 0 0 nvram_addr[1]
flabel metal2 307790 146738 307846 146794 8 FreeSans 480 90 0 0 nvram_addr[0]
flabel metal2 296954 146738 297010 146794 8 FreeSans 480 90 0 0 nvram_clk
flabel metal2 297458 146738 297514 146794 8 FreeSans 480 90 0 0 nvram_ena
flabel metal2 296450 146738 296506 146794 8 FreeSans 480 90 0 0 nvram_hr
flabel metal2 296702 146738 296758 146794 8 FreeSans 480 90 0 0 nvram_hs
flabel metal2 295946 146738 296002 146794 8 FreeSans 480 90 0 0 nvram_mem_all
flabel metal2 296198 146738 296254 146794 8 FreeSans 480 90 0 0 nvram_mem_sel
flabel metal2 315854 146738 315910 146794 8 FreeSans 480 90 0 0 nvram_rdata[31]
flabel metal2 315602 146738 315658 146794 8 FreeSans 480 90 0 0 nvram_rdata[30]
flabel metal2 315350 146738 315406 146794 8 FreeSans 480 90 0 0 nvram_rdata[29]
flabel metal2 315098 146738 315154 146794 8 FreeSans 480 90 0 0 nvram_rdata[28]
flabel metal2 314846 146738 314902 146794 8 FreeSans 480 90 0 0 nvram_rdata[27]
flabel metal2 314594 146738 314650 146794 8 FreeSans 480 90 0 0 nvram_rdata[26]
flabel metal2 314090 146738 314146 146794 8 FreeSans 480 90 0 0 nvram_rdata[24]
flabel metal2 313838 146738 313894 146794 8 FreeSans 480 90 0 0 nvram_rdata[23]
flabel metal2 313586 146738 313642 146794 8 FreeSans 480 90 0 0 nvram_rdata[22]
flabel metal2 313334 146738 313390 146794 8 FreeSans 480 90 0 0 nvram_rdata[21]
flabel metal2 313082 146738 313138 146794 8 FreeSans 480 90 0 0 nvram_rdata[20]
flabel metal2 312830 146738 312886 146794 8 FreeSans 480 90 0 0 nvram_rdata[19]
flabel metal2 312578 146738 312634 146794 8 FreeSans 480 90 0 0 nvram_rdata[18]
flabel metal2 312326 146738 312382 146794 8 FreeSans 480 90 0 0 nvram_rdata[17]
flabel metal2 312074 146738 312130 146794 8 FreeSans 480 90 0 0 nvram_rdata[16]
flabel metal2 311822 146738 311878 146794 8 FreeSans 480 90 0 0 nvram_rdata[15]
flabel metal2 311570 146738 311626 146794 8 FreeSans 480 90 0 0 nvram_rdata[14]
flabel metal2 311318 146738 311374 146794 8 FreeSans 480 90 0 0 nvram_rdata[13]
flabel metal2 311066 146738 311122 146794 8 FreeSans 480 90 0 0 nvram_rdata[12]
flabel metal2 310814 146738 310870 146794 8 FreeSans 480 90 0 0 nvram_rdata[11]
flabel metal2 310562 146738 310618 146794 8 FreeSans 480 90 0 0 nvram_rdata[10]
flabel metal2 310310 146738 310366 146794 8 FreeSans 480 90 0 0 nvram_rdata[9]
flabel metal2 310058 146738 310114 146794 8 FreeSans 480 90 0 0 nvram_rdata[8]
flabel metal2 309806 146738 309862 146794 8 FreeSans 480 90 0 0 nvram_rdata[7]
flabel metal2 309554 146738 309610 146794 8 FreeSans 480 90 0 0 nvram_rdata[6]
flabel metal2 309302 146738 309358 146794 8 FreeSans 480 90 0 0 nvram_rdata[5]
flabel metal2 309050 146738 309106 146794 8 FreeSans 480 90 0 0 nvram_rdata[4]
flabel metal2 308798 146738 308854 146794 8 FreeSans 480 90 0 0 nvram_rdata[3]
flabel metal2 308546 146738 308602 146794 8 FreeSans 480 90 0 0 nvram_rdata[2]
flabel metal2 308294 146738 308350 146794 8 FreeSans 480 90 0 0 nvram_rdata[1]
flabel metal2 308042 146738 308098 146794 8 FreeSans 480 90 0 0 nvram_rdata[0]
flabel metal2 297710 146738 297766 146794 8 FreeSans 480 90 0 0 nvram_rdy
flabel metal2 305774 146738 305830 146794 8 FreeSans 480 90 0 0 nvram_wdata[31]
flabel metal2 305522 146738 305578 146794 8 FreeSans 480 90 0 0 nvram_wdata[30]
flabel metal2 305270 146738 305326 146794 8 FreeSans 480 90 0 0 nvram_wdata[29]
flabel metal2 305018 146738 305074 146794 8 FreeSans 480 90 0 0 nvram_wdata[28]
flabel metal2 304766 146738 304822 146794 8 FreeSans 480 90 0 0 nvram_wdata[27]
flabel metal2 304514 146738 304570 146794 8 FreeSans 480 90 0 0 nvram_wdata[26]
flabel metal2 304262 146738 304318 146794 8 FreeSans 480 90 0 0 nvram_wdata[25]
flabel metal2 304010 146738 304066 146794 8 FreeSans 480 90 0 0 nvram_wdata[24]
flabel metal2 303758 146738 303814 146794 8 FreeSans 480 90 0 0 nvram_wdata[23]
flabel metal2 303506 146738 303562 146794 8 FreeSans 480 90 0 0 nvram_wdata[22]
flabel metal2 303254 146738 303310 146794 8 FreeSans 480 90 0 0 nvram_wdata[21]
flabel metal2 303002 146738 303058 146794 8 FreeSans 480 90 0 0 nvram_wdata[20]
flabel metal2 302750 146738 302806 146794 8 FreeSans 480 90 0 0 nvram_wdata[19]
flabel metal2 302498 146738 302554 146794 8 FreeSans 480 90 0 0 nvram_wdata[18]
flabel metal2 302246 146738 302302 146794 8 FreeSans 480 90 0 0 nvram_wdata[17]
flabel metal2 301994 146738 302050 146794 8 FreeSans 480 90 0 0 nvram_wdata[16]
flabel metal2 301742 146738 301798 146794 8 FreeSans 480 90 0 0 nvram_wdata[15]
flabel metal2 301490 146738 301546 146794 8 FreeSans 480 90 0 0 nvram_wdata[14]
flabel metal2 301238 146738 301294 146794 8 FreeSans 480 90 0 0 nvram_wdata[13]
flabel metal2 300986 146738 301042 146794 8 FreeSans 480 90 0 0 nvram_wdata[12]
flabel metal2 300734 146738 300790 146794 8 FreeSans 480 90 0 0 nvram_wdata[11]
flabel metal2 300482 146738 300538 146794 8 FreeSans 480 90 0 0 nvram_wdata[10]
flabel metal2 300230 146738 300286 146794 8 FreeSans 480 90 0 0 nvram_wdata[9]
flabel metal2 299978 146738 300034 146794 8 FreeSans 480 90 0 0 nvram_wdata[8]
flabel metal2 299726 146738 299782 146794 8 FreeSans 480 90 0 0 nvram_wdata[7]
flabel metal2 299474 146738 299530 146794 8 FreeSans 480 90 0 0 nvram_wdata[6]
flabel metal2 299222 146738 299278 146794 8 FreeSans 480 90 0 0 nvram_wdata[5]
flabel metal2 298970 146738 299026 146794 8 FreeSans 480 90 0 0 nvram_wdata[4]
flabel metal2 298718 146738 298774 146794 8 FreeSans 480 90 0 0 nvram_wdata[3]
flabel metal2 298466 146738 298522 146794 8 FreeSans 480 90 0 0 nvram_wdata[2]
flabel metal2 298214 146738 298270 146794 8 FreeSans 480 90 0 0 nvram_wdata[1]
flabel metal2 297962 146738 298018 146794 8 FreeSans 480 90 0 0 nvram_wdata[0]
flabel metal2 297206 146738 297262 146794 8 FreeSans 480 90 0 0 nvram_wen
flabel metal2 295694 146738 295750 146794 8 FreeSans 480 90 0 0 pass_thru
flabel metal2 233610 148120 233666 148176 8 FreeSans 480 90 0 0 flash_io2_oeb
flabel metal2 214172 148324 214228 148380 8 FreeSans 480 90 0 0 flash_io3_oeb
flabel metal2 61712 148960 61712 148960 0 FreeSans 640 90 0 0 SCK_core_lv
flabel metal3 85652 257880 85708 257936 4 FreeSans 480 0 0 0 gpio_outenb[12]
flabel metal3 90594 360266 90594 360266 0 FreeSans 480 0 0 0 gpio_in[11]
flabel metal3 85686 266582 85742 266638 4 FreeSans 480 0 0 0 gpio_outenb[0]
flabel metal3 85686 198628 85742 198684 4 FreeSans 480 0 0 0 pass_thru_csb
flabel metal3 85686 198384 85742 198440 4 FreeSans 480 0 0 0 pass_thru_sck
flabel metal3 85686 198140 85742 198196 4 FreeSans 480 0 0 0 pass_thru_sdi
flabel metal3 85686 197286 85742 197342 4 FreeSans 480 0 0 0 pass_thru_sdo
rlabel metal3 60102 128884 60158 128940 6 reg_ena
rlabel metal3 60102 129780 60158 129836 6 pll_bypass
rlabel metal3 60102 131572 60158 131628 6 pll_bias_ena
rlabel metal3 59780 136052 59836 136108 6 pll_cp_ena
rlabel metal3 59780 136276 59836 136332 6 pll_vco_ena
rlabel metal3 59780 137060 59836 137116 6 pll_vco_in
rlabel metal3 59780 137284 59836 137340 6 xtal_ena
rlabel metal3 59780 137508 59836 137564 6 prod_id[0]
rlabel metal3 59780 137732 59836 137788 6 prod_id[1]
rlabel metal3 59780 137956 59836 138012 6 prod_id[2]
rlabel metal3 59780 138180 59836 138236 6 prod_id[3]
rlabel metal3 59780 138404 59836 138460 6 prod_id[4]
rlabel metal3 59780 138628 59836 138684 6 prod_id[5]
rlabel metal3 59780 138852 59836 138908 6 prod_id[6]
rlabel metal3 59780 139076 59836 139132 6 prod_id[7]
rlabel metal3 59780 140196 59836 140252 6 mfgr_id[11]
rlabel metal3 59780 140420 59836 140476 6 mfgr_id[10]
rlabel metal3 59780 140644 59836 140700 6 mfgr_id[9]
rlabel metal3 59780 140868 59836 140924 6 mfgr_id[8]
rlabel metal3 59780 141092 59836 141148 6 mfgr_id[7]
rlabel metal3 59780 141316 59836 141372 6 mfgr_id[6]
rlabel metal3 59780 141540 59836 141596 6 mfgr_id[5]
rlabel metal3 59780 141764 59836 141820 6 mfgr_id[4]
rlabel metal3 59780 141988 59836 142044 6 mfgr_id[3]
rlabel metal3 59780 142212 59836 142268 6 mfgr_id[2]
rlabel metal3 59780 142436 59836 142492 6 mfgr_id[1]
rlabel metal3 59780 142660 59836 142716 6 mfgr_id[0]
rlabel metal3 59780 142884 59836 142940 6 mask_rev[3]
rlabel metal3 59780 143108 59836 143164 6 mask_rev[2]
rlabel metal3 59780 143332 59836 143388 6 mask_rev[1]
rlabel metal3 59780 143556 59836 143612 6 mask_rev[0]
rlabel metal3 32662 142436 32718 142492 4 sdo_enb
rlabel metal3 32662 143556 32718 143612 4 RST
flabel metal3 328706 328396 328762 328452 3 FreeSans 480 0 0 0 ram_wenb[0]
flabel metal3 328706 328152 328762 328208 3 FreeSans 480 0 0 0 ram_wenb[1]
flabel metal3 328706 327908 328762 327964 3 FreeSans 480 0 0 0 ram_wenb[2]
flabel metal3 328706 327664 328762 327720 3 FreeSans 480 0 0 0 ram_wenb[3]
flabel metal3 328706 336204 328762 336260 3 FreeSans 480 0 0 0 ram_wdata[0]
flabel metal3 328706 335960 328762 336016 3 FreeSans 480 0 0 0 ram_wdata[1]
flabel metal3 328706 335716 328762 335772 3 FreeSans 480 0 0 0 ram_wdata[2]
flabel metal3 328706 335472 328762 335528 3 FreeSans 480 0 0 0 ram_wdata[3]
flabel metal3 328706 335228 328762 335284 3 FreeSans 480 0 0 0 ram_wdata[4]
flabel metal3 328706 334984 328762 335040 3 FreeSans 480 0 0 0 ram_wdata[5]
flabel metal3 328706 334740 328762 334796 3 FreeSans 480 0 0 0 ram_wdata[6]
flabel metal3 328706 334496 328762 334552 3 FreeSans 480 0 0 0 ram_wdata[7]
flabel metal3 328706 334252 328762 334308 3 FreeSans 480 0 0 0 ram_wdata[8]
flabel metal3 328706 334008 328762 334064 3 FreeSans 480 0 0 0 ram_wdata[9]
flabel metal3 328706 333764 328762 333820 3 FreeSans 480 0 0 0 ram_wdata[10]
flabel metal3 328706 333520 328762 333576 3 FreeSans 480 0 0 0 ram_wdata[11]
flabel metal3 328706 333276 328762 333332 3 FreeSans 480 0 0 0 ram_wdata[12]
flabel metal3 328706 333032 328762 333088 3 FreeSans 480 0 0 0 ram_wdata[13]
flabel metal3 328706 332788 328762 332844 3 FreeSans 480 0 0 0 ram_wdata[14]
flabel metal3 328706 332544 328762 332600 3 FreeSans 480 0 0 0 ram_wdata[15]
flabel metal3 328706 332300 328762 332356 3 FreeSans 480 0 0 0 ram_wdata[16]
flabel metal3 328706 332056 328762 332112 3 FreeSans 480 0 0 0 ram_wdata[17]
flabel metal3 328706 331812 328762 331868 3 FreeSans 480 0 0 0 ram_wdata[18]
flabel metal3 328706 331568 328762 331624 3 FreeSans 480 0 0 0 ram_wdata[19]
flabel metal3 328706 331324 328762 331380 3 FreeSans 480 0 0 0 ram_wdata[20]
flabel metal3 328706 331080 328762 331136 3 FreeSans 480 0 0 0 ram_wdata[21]
flabel metal3 328706 330836 328762 330892 3 FreeSans 480 0 0 0 ram_wdata[22]
flabel metal3 328706 330592 328762 330648 3 FreeSans 480 0 0 0 ram_wdata[23]
flabel metal3 328706 330348 328762 330404 3 FreeSans 480 0 0 0 ram_wdata[24]
flabel metal3 328706 330104 328762 330160 3 FreeSans 480 0 0 0 ram_wdata[25]
flabel metal3 328706 329860 328762 329916 3 FreeSans 480 0 0 0 ram_wdata[26]
flabel metal3 328706 329616 328762 329672 3 FreeSans 480 0 0 0 ram_wdata[27]
flabel metal3 328706 329372 328762 329428 3 FreeSans 480 0 0 0 ram_wdata[28]
flabel metal3 328706 329128 328762 329184 3 FreeSans 480 0 0 0 ram_wdata[29]
flabel metal3 328706 328884 328762 328940 3 FreeSans 480 0 0 0 ram_wdata[30]
flabel metal3 328706 328640 328762 328696 3 FreeSans 480 0 0 0 ram_wdata[31]
flabel metal3 328706 316928 328762 316984 3 FreeSans 480 0 0 0 ram_rdata[0]
flabel metal3 328706 317172 328762 317228 3 FreeSans 480 0 0 0 ram_rdata[1]
flabel metal3 328706 317416 328762 317472 3 FreeSans 480 0 0 0 ram_rdata[2]
flabel metal3 328706 317660 328762 317716 3 FreeSans 480 0 0 0 ram_rdata[3]
flabel metal3 328706 317904 328762 317960 3 FreeSans 480 0 0 0 ram_rdata[4]
flabel metal3 328706 318148 328762 318204 3 FreeSans 480 0 0 0 ram_rdata[5]
flabel metal3 328706 318392 328762 318448 3 FreeSans 480 0 0 0 ram_rdata[6]
flabel metal3 328706 318636 328762 318692 3 FreeSans 480 0 0 0 ram_rdata[7]
flabel metal3 328706 318880 328762 318936 3 FreeSans 480 0 0 0 ram_rdata[8]
flabel metal3 328706 319124 328762 319180 3 FreeSans 480 0 0 0 ram_rdata[9]
flabel metal3 328706 319368 328762 319424 3 FreeSans 480 0 0 0 ram_rdata[10]
flabel metal3 328706 319612 328762 319668 3 FreeSans 480 0 0 0 ram_rdata[11]
flabel metal3 328706 319856 328762 319912 3 FreeSans 480 0 0 0 ram_rdata[12]
flabel metal3 328706 320100 328762 320156 3 FreeSans 480 0 0 0 ram_rdata[13]
flabel metal3 328706 320344 328762 320400 3 FreeSans 480 0 0 0 ram_rdata[14]
flabel metal3 328706 320588 328762 320644 3 FreeSans 480 0 0 0 ram_rdata[15]
flabel metal3 328706 320832 328762 320888 3 FreeSans 480 0 0 0 ram_rdata[16]
flabel metal3 328706 321076 328762 321132 3 FreeSans 480 0 0 0 ram_rdata[17]
flabel metal3 328706 321320 328762 321376 3 FreeSans 480 0 0 0 ram_rdata[18]
flabel metal3 328706 321564 328762 321620 3 FreeSans 480 0 0 0 ram_rdata[19]
flabel metal3 328706 321808 328762 321864 3 FreeSans 480 0 0 0 ram_rdata[20]
flabel metal3 328706 322052 328762 322108 3 FreeSans 480 0 0 0 ram_rdata[21]
flabel metal3 328706 322296 328762 322352 3 FreeSans 480 0 0 0 ram_rdata[22]
flabel metal3 328706 322540 328762 322596 3 FreeSans 480 0 0 0 ram_rdata[23]
flabel metal3 328706 322784 328762 322840 3 FreeSans 480 0 0 0 ram_rdata[24]
flabel metal3 328706 323028 328762 323084 3 FreeSans 480 0 0 0 ram_rdata[25]
flabel metal3 328706 323272 328762 323328 3 FreeSans 480 0 0 0 ram_rdata[26]
flabel metal3 328706 323516 328762 323572 3 FreeSans 480 0 0 0 ram_rdata[27]
flabel metal3 328706 323760 328762 323816 3 FreeSans 480 0 0 0 ram_rdata[28]
flabel metal3 328706 324004 328762 324060 3 FreeSans 480 0 0 0 ram_rdata[29]
flabel metal3 328706 324248 328762 324304 3 FreeSans 480 0 0 0 ram_rdata[30]
flabel metal3 328706 324492 328762 324548 3 FreeSans 480 0 0 0 ram_rdata[31]
flabel metal3 328706 327420 328762 327476 3 FreeSans 480 0 0 0 ram_addr[0]
flabel metal3 328706 327176 328762 327232 3 FreeSans 480 0 0 0 ram_addr[1]
flabel metal3 328706 326932 328762 326988 3 FreeSans 480 0 0 0 ram_addr[2]
flabel metal3 328706 326688 328762 326744 3 FreeSans 480 0 0 0 ram_addr[3]
flabel metal3 328706 326444 328762 326500 3 FreeSans 480 0 0 0 ram_addr[4]
flabel metal3 328706 326200 328762 326256 3 FreeSans 480 0 0 0 ram_addr[5]
flabel metal3 328706 325956 328762 326012 3 FreeSans 480 0 0 0 ram_addr[6]
flabel metal3 328706 325712 328762 325768 3 FreeSans 480 0 0 0 ram_addr[7]
flabel metal3 328706 325468 328762 325524 3 FreeSans 480 0 0 0 ram_addr[8]
flabel metal3 328706 325224 328762 325280 3 FreeSans 480 0 0 0 ram_addr[9]
flabel metal3 328706 324980 328762 325036 3 FreeSans 480 0 0 0 ram_addr[10]
flabel metal3 328706 324736 328762 324792 3 FreeSans 480 0 0 0 ram_addr[11]
flabel metal3 85652 245436 85708 245492 4 FreeSans 480 0 0 0 gpio_out[15]
flabel metal3 85652 245680 85708 245736 4 FreeSans 480 0 0 0 gpio_out[14]
flabel metal3 85652 245924 85708 245980 4 FreeSans 480 0 0 0 gpio_out[13]
flabel metal3 85652 246168 85708 246224 4 FreeSans 480 0 0 0 gpio_out[12]
flabel metal3 85652 246412 85708 246468 4 FreeSans 480 0 0 0 gpio_out[11]
flabel metal3 85652 246656 85708 246712 4 FreeSans 480 0 0 0 gpio_out[10]
flabel metal3 85652 246900 85708 246956 4 FreeSans 480 0 0 0 gpio_out[9]
flabel metal3 85652 247144 85708 247200 4 FreeSans 480 0 0 0 gpio_out[8]
flabel metal3 85652 247388 85708 247444 4 FreeSans 480 0 0 0 gpio_out[7]
flabel metal3 85652 247632 85708 247688 4 FreeSans 480 0 0 0 gpio_out[6]
flabel metal3 85652 247876 85708 247932 4 FreeSans 480 0 0 0 gpio_out[5]
flabel metal3 85652 248120 85708 248176 4 FreeSans 480 0 0 0 gpio_out[4]
flabel metal3 85652 248364 85708 248420 4 FreeSans 480 0 0 0 gpio_out[3]
flabel metal3 85652 248608 85708 248664 4 FreeSans 480 0 0 0 gpio_out[2]
flabel metal3 85652 248852 85708 248908 4 FreeSans 480 0 0 0 gpio_out[1]
flabel metal3 85652 249096 85708 249152 4 FreeSans 480 0 0 0 gpio_out[0]
flabel metal3 85652 257148 85708 257204 4 FreeSans 480 0 0 0 gpio_outenb[15]
flabel metal3 85652 257392 85708 257448 4 FreeSans 480 0 0 0 gpio_outenb[14]
flabel metal3 85652 257636 85708 257692 4 FreeSans 480 0 0 0 gpio_outenb[13]
flabel metal3 85652 258124 85708 258180 4 FreeSans 480 0 0 0 gpio_outenb[11]
flabel metal3 85652 258368 85708 258424 4 FreeSans 480 0 0 0 gpio_outenb[10]
flabel metal3 85652 258612 85708 258668 4 FreeSans 480 0 0 0 gpio_outenb[9]
flabel metal3 85652 258856 85708 258912 4 FreeSans 480 0 0 0 gpio_outenb[8]
flabel metal3 85652 259100 85708 259156 4 FreeSans 480 0 0 0 gpio_outenb[7]
flabel metal3 85652 259344 85708 259400 4 FreeSans 480 0 0 0 gpio_outenb[6]
flabel metal3 85652 259588 85708 259644 4 FreeSans 480 0 0 0 gpio_outenb[5]
flabel metal3 85652 259832 85708 259888 4 FreeSans 480 0 0 0 gpio_outenb[4]
flabel metal3 85652 260076 85708 260132 4 FreeSans 480 0 0 0 gpio_outenb[3]
flabel metal3 85652 260320 85708 260376 4 FreeSans 480 0 0 0 gpio_outenb[2]
flabel metal3 85652 260564 85708 260620 4 FreeSans 480 0 0 0 gpio_outenb[1]
flabel metal3 85652 249340 85708 249396 4 FreeSans 480 0 0 0 gpio_pulldownb[15]
flabel metal3 85652 249584 85708 249640 4 FreeSans 480 0 0 0 gpio_pulldownb[14]
flabel metal3 85652 249828 85708 249884 4 FreeSans 480 0 0 0 gpio_pulldownb[13]
flabel metal3 85652 250072 85708 250128 4 FreeSans 480 0 0 0 gpio_pulldownb[12]
flabel metal3 85652 250316 85708 250372 4 FreeSans 480 0 0 0 gpio_pulldownb[11]
flabel metal3 85652 250560 85708 250616 4 FreeSans 480 0 0 0 gpio_pulldownb[10]
flabel metal3 85652 250804 85708 250860 4 FreeSans 480 0 0 0 gpio_pulldownb[9]
flabel metal3 85652 251048 85708 251104 4 FreeSans 480 0 0 0 gpio_pulldownb[8]
flabel metal3 85652 251292 85708 251348 4 FreeSans 480 0 0 0 gpio_pulldownb[7]
flabel metal3 85652 251536 85708 251592 4 FreeSans 480 0 0 0 gpio_pulldownb[6]
flabel metal3 85652 251780 85708 251836 4 FreeSans 480 0 0 0 gpio_pulldownb[5]
flabel metal3 85652 252024 85708 252080 4 FreeSans 480 0 0 0 gpio_pulldownb[4]
flabel metal3 85652 252268 85708 252324 4 FreeSans 480 0 0 0 gpio_pulldownb[3]
flabel metal3 85652 252512 85708 252568 4 FreeSans 480 0 0 0 gpio_pulldownb[2]
flabel metal3 85652 252756 85708 252812 4 FreeSans 480 0 0 0 gpio_pulldownb[1]
flabel metal3 85652 253000 85708 253056 4 FreeSans 480 0 0 0 gpio_pulldownb[0]
flabel metal3 85652 256904 85708 256960 4 FreeSans 480 0 0 0 gpio_pullupb[15]
flabel metal3 85652 256660 85708 256716 4 FreeSans 480 0 0 0 gpio_pullupb[14]
flabel metal3 85652 256416 85708 256472 4 FreeSans 480 0 0 0 gpio_pullupb[13]
flabel metal3 85652 256172 85708 256228 4 FreeSans 480 0 0 0 gpio_pullupb[12]
flabel metal3 85652 255928 85708 255984 4 FreeSans 480 0 0 0 gpio_pullupb[11]
flabel metal3 85652 255684 85708 255740 4 FreeSans 480 0 0 0 gpio_pullupb[10]
flabel metal3 85652 255440 85708 255496 4 FreeSans 480 0 0 0 gpio_pullupb[9]
flabel metal3 85652 255196 85708 255252 4 FreeSans 480 0 0 0 gpio_pullupb[8]
flabel metal3 85652 254952 85708 255008 4 FreeSans 480 0 0 0 gpio_pullupb[7]
flabel metal3 85652 254708 85708 254764 4 FreeSans 480 0 0 0 gpio_pullupb[6]
flabel metal3 85652 254464 85708 254520 4 FreeSans 480 0 0 0 gpio_pullupb[5]
flabel metal3 85652 254220 85708 254276 4 FreeSans 480 0 0 0 gpio_pullupb[4]
flabel metal3 85652 253976 85708 254032 4 FreeSans 480 0 0 0 gpio_pullupb[3]
flabel metal3 85652 253732 85708 253788 4 FreeSans 480 0 0 0 gpio_pullupb[2]
flabel metal3 85652 253488 85708 253544 4 FreeSans 480 0 0 0 gpio_pullupb[1]
flabel metal3 85652 253244 85708 253300 4 FreeSans 480 0 0 0 gpio_pullupb[0]
flabel metal3 85652 351210 85708 351266 4 FreeSans 480 0 0 0 adc0_data[9]
flabel metal3 85652 350966 85708 351022 4 FreeSans 480 0 0 0 adc0_data[8]
flabel metal3 85652 350722 85708 350778 4 FreeSans 480 0 0 0 adc0_data[7]
flabel metal3 85652 350478 85708 350534 4 FreeSans 480 0 0 0 adc0_data[6]
flabel metal3 85652 350234 85708 350290 4 FreeSans 480 0 0 0 adc0_data[5]
flabel metal3 85652 349990 85708 350046 4 FreeSans 480 0 0 0 adc0_data[4]
flabel metal3 85652 349746 85708 349802 4 FreeSans 480 0 0 0 adc0_data[3]
flabel metal3 85652 349502 85708 349558 4 FreeSans 480 0 0 0 adc0_data[2]
flabel metal3 85652 349258 85708 349314 4 FreeSans 480 0 0 0 adc0_data[1]
flabel metal3 85652 349014 85708 349070 4 FreeSans 480 0 0 0 adc0_data[0]
flabel metal3 85652 356822 85708 356878 4 FreeSans 480 0 0 0 adc0_inputsrc[1]
flabel metal3 85652 357066 85708 357122 4 FreeSans 480 0 0 0 adc0_inputsrc[0]
flabel metal3 85652 351698 85708 351754 4 FreeSans 480 0 0 0 adc1_data[8]
flabel metal3 85652 351942 85708 351998 4 FreeSans 480 0 0 0 adc1_data[7]
flabel metal3 85652 352186 85708 352242 4 FreeSans 480 0 0 0 adc1_data[6]
flabel metal3 85652 352430 85708 352486 4 FreeSans 480 0 0 0 adc1_data[5]
flabel metal3 85652 352674 85708 352730 4 FreeSans 480 0 0 0 adc1_data[4]
flabel metal3 85652 352918 85708 352974 4 FreeSans 480 0 0 0 adc1_data[3]
flabel metal3 85652 353162 85708 353218 4 FreeSans 480 0 0 0 adc1_data[2]
flabel metal3 85652 353406 85708 353462 4 FreeSans 480 0 0 0 adc1_data[1]
flabel metal3 85652 353650 85708 353706 4 FreeSans 480 0 0 0 adc1_data[0]
flabel metal3 85652 356578 85708 356634 4 FreeSans 480 0 0 0 adc1_inputsrc[1]
flabel metal3 85652 356334 85708 356390 4 FreeSans 480 0 0 0 adc1_inputsrc[0]
flabel metal3 85652 356090 85708 356146 4 FreeSans 480 0 0 0 dac_value[9]
flabel metal3 85652 355846 85708 355902 4 FreeSans 480 0 0 0 dac_value[8]
flabel metal3 85652 355602 85708 355658 4 FreeSans 480 0 0 0 dac_value[7]
flabel metal3 85652 355358 85708 355414 4 FreeSans 480 0 0 0 dac_value[6]
flabel metal3 85652 355114 85708 355170 4 FreeSans 480 0 0 0 dac_value[5]
flabel metal3 85652 354870 85708 354926 4 FreeSans 480 0 0 0 dac_value[4]
flabel metal3 85652 354626 85708 354682 4 FreeSans 480 0 0 0 dac_value[3]
flabel metal3 85652 354382 85708 354438 4 FreeSans 480 0 0 0 dac_value[2]
flabel metal3 85652 354138 85708 354194 4 FreeSans 480 0 0 0 dac_value[1]
flabel metal3 85652 353894 85708 353950 4 FreeSans 480 0 0 0 dac_value[0]
flabel metal3 85652 348770 85708 348826 4 FreeSans 480 0 0 0 ext_reset
flabel metal3 85652 348282 85708 348338 4 FreeSans 480 0 0 0 irq_pin
flabel metal3 85652 317782 85708 317838 4 FreeSans 480 0 0 0 irq_spi
flabel metal3 85652 348526 85708 348582 4 FreeSans 480 0 0 0 reset
flabel metal3 85652 314854 85708 314910 4 FreeSans 480 0 0 0 spi_ro_config[7]
flabel metal3 85652 315098 85708 315154 4 FreeSans 480 0 0 0 spi_ro_config[6]
flabel metal3 85652 315342 85708 315398 4 FreeSans 480 0 0 0 spi_ro_config[5]
flabel metal3 85652 315586 85708 315642 4 FreeSans 480 0 0 0 spi_ro_config[4]
flabel metal3 85652 315830 85708 315886 4 FreeSans 480 0 0 0 spi_ro_config[3]
flabel metal3 85652 316074 85708 316130 4 FreeSans 480 0 0 0 spi_ro_config[2]
flabel metal3 85652 316806 85708 316862 4 FreeSans 480 0 0 0 spi_ro_mask_rev[3]
flabel metal3 85652 317050 85708 317106 4 FreeSans 480 0 0 0 spi_ro_mask_rev[2]
flabel metal3 85652 317294 85708 317350 4 FreeSans 480 0 0 0 spi_ro_mask_rev[1]
flabel metal3 85652 346818 85708 346874 4 FreeSans 480 0 0 0 spi_ro_pll_bias_ena
flabel metal3 85652 347306 85708 347362 4 FreeSans 480 0 0 0 spi_ro_pll_cp_ena
flabel metal3 85652 347062 85708 347118 4 FreeSans 480 0 0 0 spi_ro_pll_vco_ena
flabel metal3 85652 305582 85708 305638 4 FreeSans 480 0 0 0 spi_ro_prod_id[7]
flabel metal3 85652 313146 85708 313202 4 FreeSans 480 0 0 0 spi_ro_prod_id[6]
flabel metal3 85652 313390 85708 313446 4 FreeSans 480 0 0 0 spi_ro_prod_id[5]
flabel metal3 85652 313634 85708 313690 4 FreeSans 480 0 0 0 spi_ro_prod_id[4]
flabel metal3 85652 313878 85708 313934 4 FreeSans 480 0 0 0 spi_ro_prod_id[3]
flabel metal3 85652 314122 85708 314178 4 FreeSans 480 0 0 0 spi_ro_prod_id[2]
flabel metal3 85652 314366 85708 314422 4 FreeSans 480 0 0 0 spi_ro_prod_id[1]
flabel metal3 85652 347550 85708 347606 4 FreeSans 480 0 0 0 spi_ro_reg_ena
flabel metal3 85652 347794 85708 347850 4 FreeSans 480 0 0 0 spi_ro_xtal_ena
flabel metal3 85652 348038 85708 348094 4 FreeSans 480 0 0 0 trap
flabel metal3 90594 359778 90594 359778 0 FreeSans 480 0 0 0 gpio_in[9]
flabel metal3 90594 360022 90594 360022 0 FreeSans 480 0 0 0 gpio_in[10]
flabel metal3 90594 360510 90594 360510 0 FreeSans 480 0 0 0 gpio_in[12]
flabel metal3 90594 360754 90594 360754 0 FreeSans 480 0 0 0 gpio_in[13]
flabel metal3 90594 360998 90594 360998 0 FreeSans 480 0 0 0 gpio_in[14]
flabel metal3 90594 361242 90594 361242 0 FreeSans 480 0 0 0 gpio_in[15]
flabel metal3 90594 361486 90594 361486 0 FreeSans 480 0 0 0 adc0_done
flabel metal3 90594 361730 90594 361730 0 FreeSans 480 0 0 0 adc1_done
flabel metal3 90594 362218 90594 362218 0 FreeSans 480 0 0 0 rosc_in
flabel metal3 90594 362462 90594 362462 0 FreeSans 480 0 0 0 comp_in
flabel metal3 90594 362706 90594 362706 0 FreeSans 480 0 0 0 adc0_ena
flabel metal3 90594 362950 90594 362950 0 FreeSans 480 0 0 0 adc0_convert
flabel metal3 90594 363194 90594 363194 0 FreeSans 480 0 0 0 adc0_clk
flabel metal3 90594 363438 90594 363438 0 FreeSans 480 0 0 0 adc1_ena
flabel metal3 90594 363682 90594 363682 0 FreeSans 480 0 0 0 adc1_convert
flabel metal3 90594 363926 90594 363926 0 FreeSans 480 0 0 0 adc1_clk
flabel metal3 90594 364170 90594 364170 0 FreeSans 480 0 0 0 dac_ena
flabel metal3 90594 364414 90594 364414 0 FreeSans 480 0 0 0 analog_out_sel
flabel metal3 90594 364658 90594 364658 0 FreeSans 480 0 0 0 opamp_ena
flabel metal3 90594 364902 90594 364902 0 FreeSans 480 0 0 0 opamp_bias_ena
flabel metal3 90594 365146 90594 365146 0 FreeSans 480 0 0 0 bg_ena
flabel metal3 90594 365390 90594 365390 0 FreeSans 480 0 0 0 comp_ena
flabel metal3 90594 365634 90594 365634 0 FreeSans 480 0 0 0 rcosc_ena
flabel metal3 90594 366122 90594 366122 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[11]
flabel metal3 90594 366366 90594 366366 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[10]
flabel metal3 90594 366610 90594 366610 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[9]
flabel metal3 90594 366854 90594 366854 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[8]
flabel metal3 90594 367098 90594 367098 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[7]
flabel metal3 90594 367342 90594 367342 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[6]
flabel metal3 90594 367586 90594 367586 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[5]
flabel metal3 90594 367830 90594 367830 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[4]
flabel metal3 90594 368074 90594 368074 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[3]
flabel metal3 90594 368318 90594 368318 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[2]
flabel metal3 90594 368562 90594 368562 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[1]
flabel metal3 90594 368806 90594 368806 0 FreeSans 480 0 0 0 spi_ro_mfgr_id[0]
flabel metal3 90594 369050 90594 369050 0 FreeSans 480 0 0 0 comp_pinputsrc[1]
flabel metal3 90594 369294 90594 369294 0 FreeSans 480 0 0 0 comp_pinputsrc[0]
flabel metal3 90594 369538 90594 369538 0 FreeSans 480 0 0 0 spi_ro_pll_trim[0]
flabel metal3 90594 369782 90594 369782 0 FreeSans 480 0 0 0 spi_ro_pll_trim[1]
flabel metal3 90594 370026 90594 370026 0 FreeSans 480 0 0 0 spi_ro_pll_trim[2]
flabel metal3 90594 370270 90594 370270 0 FreeSans 480 0 0 0 spi_ro_pll_trim[3]
flabel metal3 90594 370514 90594 370514 0 FreeSans 480 0 0 0 comp_ninputsrc[0]
flabel metal3 90594 370758 90594 370758 0 FreeSans 480 0 0 0 comp_ninputsrc[1]
flabel metal3 85652 314610 85708 314666 4 FreeSans 480 0 0 0 spi_ro_prod_id[0]
flabel metal3 85652 317538 85708 317594 4 FreeSans 480 0 0 0 spi_ro_mask_rev[0]
flabel via2 314342 146738 314398 146794 8 FreeSans 480 90 0 0 nvram_rdata[25]
flabel metal2 81872 163856 81872 163856 0 FreeSans 640 90 0 0 adc1_clock
flabel metal2 81760 163856 81760 163856 0 FreeSans 640 90 0 0 adc1_start
flabel metal2 81648 163856 81648 163856 0 FreeSans 640 90 0 0 adc1_ena
flabel metal2 81536 163856 81536 163856 0 FreeSans 640 90 0 0 adc1_done
flabel metal2 81424 163856 81424 163856 0 FreeSans 640 90 0 0 adc1_data[0]
flabel metal2 81312 164080 81312 164080 0 FreeSans 640 90 0 0 adc1_data[1]
flabel metal2 81200 164080 81200 164080 0 FreeSans 640 90 0 0 adc1_data[2]
flabel metal2 81088 164080 81088 164080 0 FreeSans 640 90 0 0 adc1_data[3]
flabel metal2 80976 164080 80976 164080 0 FreeSans 640 90 0 0 adc1_data[4]
flabel metal2 80864 164080 80864 164080 0 FreeSans 640 90 0 0 adc1_data[5]
flabel metal2 80752 164080 80752 164080 0 FreeSans 640 90 0 0 adc1_data[6]
flabel metal2 80640 164080 80640 164080 0 FreeSans 640 90 0 0 adc1_data[7]
flabel metal2 80528 164080 80528 164080 0 FreeSans 640 90 0 0 adc1_data[8]
flabel metal2 80416 164080 80416 164080 0 FreeSans 640 90 0 0 adc1_data[9]
flabel metal2 83440 207536 83440 207536 0 FreeSans 640 90 0 0 adc0_clock
flabel metal2 83328 207536 83328 207536 0 FreeSans 640 90 0 0 adc0_start
flabel metal2 83216 207536 83216 207536 0 FreeSans 640 90 0 0 adc0_ena
flabel metal2 83104 207536 83104 207536 0 FreeSans 640 90 0 0 adc0_done
flabel metal2 82992 207536 82992 207536 0 FreeSans 640 90 0 0 adc0_data[0]
flabel metal2 82880 207536 82880 207536 0 FreeSans 640 90 0 0 adc0_data[1]
flabel metal2 82768 207536 82768 207536 0 FreeSans 640 90 0 0 adc0_data[2]
flabel metal2 82656 207536 82656 207536 0 FreeSans 640 90 0 0 adc0_data[3]
flabel metal2 82544 207536 82544 207536 0 FreeSans 640 90 0 0 adc0_data[4]
flabel metal2 82432 207536 82432 207536 0 FreeSans 640 90 0 0 adc0_data[5]
flabel metal2 82320 207536 82320 207536 0 FreeSans 640 90 0 0 adc0_data[6]
flabel metal2 82208 207536 82208 207536 0 FreeSans 640 90 0 0 adc0_data[7]
flabel metal2 82096 207536 82096 207536 0 FreeSans 640 90 0 0 adc0_data[8]
flabel metal2 81984 207536 81984 207536 0 FreeSans 640 90 0 0 adc0_data[9]
flabel metal3 85652 351454 85708 351510 4 FreeSans 480 0 0 0 adc1_data[9]
flabel metal3 101693 106823 101693 106823 0 FreeSans 800 0 0 0 bias10u
flabel metal3 101692 106522 101692 106522 0 FreeSans 800 0 0 0 bias5u
flabel metaltp 45800 369200 45800 369200 0 FreeSans 8000 0 0 0 VDD3V3
flabel metaltp 46200 362000 46200 362000 0 FreeSans 8000 0 0 0 VSS
flabel metaltpl 76986 119196 76986 119196 0 FreeSans 5040 90 0 0 VDD3V3
flabel metaltpl 84420 119070 84420 119070 0 FreeSans 5040 90 0 0 VSS
flabel metaltpl 111132 118566 111132 118566 0 FreeSans 5040 90 0 0 VDD1V8
flabel metal2 66640 132272 66640 132272 0 FreeSans 640 90 0 0 dground
flabel metal1 429296 392560 439824 405776 0 FreeSans 16000 90 0 0 VDD3V3
port 0 nsew
flabel metal1 446096 392560 456624 405776 0 FreeSans 16000 90 0 0 VSS
flabel metal1 493584 351120 506688 361648 0 FreeSans 16000 0 0 0 VSS
port 2 nsew
flabel metal1 493584 243936 506688 254464 0 FreeSans 16000 0 0 0 ser_rx
port 11 nsew
flabel metal1 493584 227136 506688 237664 0 FreeSans 16000 0 0 0 ser_tx
port 10 nsew
flabel metal1 493584 136752 506688 147280 0 FreeSans 16000 0 0 0 i2c_scl
port 13 nsew
flabel metal1 493584 119952 506688 130480 0 FreeSans 16000 0 0 0 i2c_sda
port 12 nsew
flabel metal1 493584 46368 506688 56896 0 FreeSans 16000 0 0 0 irq
port 18 nsew
flabel metal1 468944 7840 479472 20944 0 FreeSans 16000 90 0 0 XCLK
port 5 nsew
flabel metal1 418096 7840 428624 20944 0 FreeSans 16000 90 0 0 flash_io3
port 40 nsew
flabel metal1 401296 7840 411824 20944 0 FreeSans 16000 90 0 0 flash_io2
port 39 nsew
flabel metal1 384496 7840 395024 20944 0 FreeSans 16000 90 0 0 flash_io1
port 38 nsew
flabel metal1 367696 7840 378224 20944 0 FreeSans 16000 90 0 0 flash_io0
port 37 nsew
flabel metal1 330960 7840 341488 20944 0 FreeSans 16000 90 0 0 flash_csb
port 35 nsew
flabel metal1 314160 7840 324688 20944 0 FreeSans 16000 90 0 0 flash_clk
port 36 nsew
flabel metal1 287280 7840 297808 20944 0 FreeSans 16000 90 0 0 VDD1V8
port 1 nsew
flabel metaltpl 12320 65296 16464 68544 0 FreeSans 16000 0 0 0 XO
port 4 nsew
flabel metaltpl 12768 104160 16240 107184 0 FreeSans 16000 0 0 0 XI
port 3 nsew
flabel metal1 7840 117152 20944 127680 0 FreeSans 16000 0 0 0 nvref_ext
port 48 nsew
flabel metal1 7840 143920 20944 154448 0 FreeSans 16000 0 0 0 adc0_in
port 43 nsew
flabel metal1 7840 160720 20944 171248 0 FreeSans 16000 0 0 0 adc1_in
port 44 nsew
flabel metal1 7840 177520 20944 188048 0 FreeSans 16000 0 0 0 adc_low
port 42 nsew
flabel metal1 7840 194320 20944 204848 0 FreeSans 16000 0 0 0 adc_high
port 41 nsew
flabel metal1 7840 211120 20944 221648 0 FreeSans 16000 0 0 0 analog_out
port 45 nsew
flabel metal1 7840 227920 20944 238448 0 FreeSans 16000 0 0 0 comp_inn
port 47 nsew
flabel metal1 7840 244720 20944 255248 0 FreeSans 16000 0 0 0 comp_inp
port 46 nsew
flabel metal1 7840 273840 20944 284368 0 FreeSans 16000 0 0 0 gpio[15]
port 19 nsew
flabel metal1 7840 290752 20944 301280 0 FreeSans 16000 0 0 0 gpio[14]
port 20 nsew
flabel metal1 7840 307552 20944 318080 0 FreeSans 16000 0 0 0 gpio[13]
port 21 nsew
flabel metal1 7840 324352 20944 334880 0 FreeSans 16000 0 0 0 gpio[12]
port 22 nsew
flabel metal1 35168 392560 45584 405664 0 FreeSans 16000 90 0 0 gpio[11]
port 23 nsew
flabel metal1 51968 392560 62384 405664 0 FreeSans 16000 90 0 0 gpio[10]
port 24 nsew
flabel metal1 68768 392560 79184 405664 0 FreeSans 16000 90 0 0 gpio[9]
port 25 nsew
flabel metal1 85568 392560 95984 405664 0 FreeSans 16000 90 0 0 gpio[8]
port 26 nsew
flabel metal1 102368 392560 112784 405664 0 FreeSans 16000 90 0 0 gpio[7]
port 27 nsew
flabel metal1 119168 392560 129584 405664 0 FreeSans 16000 90 0 0 gpio[6]
port 28 nsew
flabel metal1 135968 392560 146384 405664 0 FreeSans 16000 90 0 0 gpio[5]
port 29 nsew
flabel metal1 192752 392560 203168 405664 0 FreeSans 16000 90 0 0 gpio[4]
port 30 nsew
flabel metal1 209552 392560 219968 405664 0 FreeSans 16000 90 0 0 gpio[3]
port 31 nsew
flabel metal1 236432 392560 246848 405664 0 FreeSans 16000 90 0 0 gpio[2]
port 32 nsew
flabel metal1 253232 392560 263648 405664 0 FreeSans 16000 90 0 0 gpio[1]
port 33 nsew
flabel metal1 269920 392560 280336 405664 0 FreeSans 16000 90 0 0 gpio[0]
port 34 nsew
flabel metal1 493584 367920 506688 378448 0 FreeSans 16000 0 0 0 spi_sdi
port 14 nsew
flabel metal1 493584 334320 506688 344848 0 FreeSans 16000 0 0 0 spi_csb
port 15 nsew
flabel metal1 493584 317520 506688 328048 0 FreeSans 16000 0 0 0 spi_sck
port 16 nsew
flabel metal1 493584 300720 506688 311248 0 FreeSans 16000 0 0 0 spi_sdo
port 17 nsew
rlabel metal3 60102 128212 60158 128268 6 spi_reset
rlabel metal3 59780 139972 59836 140028 6 spi_pass_thru_sdo
rlabel metal3 59780 139748 59836 139804 6 spi_pass_thru_sck
rlabel metal3 59780 139524 59836 139580 6 spi_pass_thru_csb
rlabel metal3 59780 139300 59836 139356 6 spi_pass_thru_sdi
rlabel metal3 32662 143332 32718 143388 4 SCK_core
rlabel metal3 32662 143108 32718 143164 4 SDI_core
rlabel metal3 32662 142884 32718 142940 4 CSB_core
rlabel metal3 32662 142660 32718 142716 4 SDO_core
flabel metal2 294182 146738 294238 146794 8 FreeSans 480 90 0 0 flash_clk_core
flabel metal2 295442 146738 295498 146794 8 FreeSans 480 90 0 0 flash_csb_core
flabel metal2 314342 359628 314398 359684 6 FreeSans 480 90 0 0 ser_rx_core
flabel metal2 314594 359628 314650 359684 6 FreeSans 480 90 0 0 ser_tx_core
rlabel metal3 60102 126196 60158 126252 6 irq_core
rlabel metal3 60102 127988 60158 128044 6 spi_trap_in
flabel metal3 85652 346574 85708 346630 4 FreeSans 480 0 0 0 spi_sck_core
flabel metaltpl 321858 369904 321858 369904 0 FreeSans 8000 90 0 0 VDD1V8
flabel metal2 85332 146159 85332 146159 0 FreeSans 640 90 0 0 reg1_enb
flabel metal2 86686 146174 86686 146174 0 FreeSans 640 90 0 0 reg1_ena
flabel metal2 68320 136528 68320 136528 0 FreeSans 640 90 0 0 spare_dg
flabel metal2 84903 146167 84903 146167 0 FreeSans 640 90 0 0 reg0_enb
flabel metal2 86004 146159 86004 146159 0 FreeSans 640 90 0 0 reg0_ena
flabel metal1 87536 7840 98064 20944 0 FreeSans 16000 90 0 0 SCK
port 9 nsew
flabel metal1 70736 7840 81264 20944 0 FreeSans 16000 90 0 0 CSB
port 8 nsew
flabel metal1 53936 7840 64464 20944 0 FreeSans 16000 90 0 0 SDI
port 6 nsew
flabel metal1 37136 7840 47664 20944 0 FreeSans 16000 90 0 0 SDO
port 7 nsew
<< end >>
