magic
tech EFXH018D
timestamp 1494891594
<< metal2 >>
tri 160 1920 480 2240 se
rect 480 2024 1648 2240
tri 480 1920 584 2024 nw
tri 1544 1920 1648 2024 ne
tri 1648 1968 1920 2240 sw
rect 1648 1920 1920 1968
tri -104 1648 160 1920 se
rect -104 1600 160 1648
tri 160 1600 480 1920 nw
tri 1648 1648 1920 1920 ne
tri 1920 1648 2240 1968 sw
rect -104 480 104 1600
tri 104 1544 160 1600 nw
rect 528 1204 632 1600
tri 632 1204 1028 1600 sw
tri 1100 1204 1496 1600 se
rect 1496 1204 1600 1600
tri 1920 1544 2024 1648 ne
rect 528 1144 1600 1204
tri 104 480 208 584 sw
rect 528 528 744 1144
tri 824 960 1008 1144 ne
rect 1008 960 1120 1144
tri 1120 960 1304 1144 nw
rect 1384 528 1600 1144
tri 1920 480 2024 584 se
rect 2024 480 2240 1648
tri -104 160 208 480 ne
tri 208 160 528 480 sw
tri 1600 160 1920 480 se
tri 1920 160 2240 480 nw
tri 208 -104 480 160 ne
rect 480 104 528 160
tri 528 104 584 160 sw
tri 1544 104 1600 160 se
rect 1600 104 1648 160
rect 480 -104 1648 104
tri 1648 -104 1920 160 nw
<< end >>
