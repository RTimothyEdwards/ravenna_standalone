magic
tech EFXH018D
timestamp 1533305873
<< mimcap >>
rect -11240 5225 -9240 5240
rect -11240 2755 -11225 5225
rect -9255 2755 -9240 5225
rect -11240 2740 -9240 2755
rect -8975 5225 -6975 5240
rect -8975 2755 -8960 5225
rect -6990 2755 -6975 5225
rect -8975 2740 -6975 2755
rect -6710 5225 -4710 5240
rect -6710 2755 -6695 5225
rect -4725 2755 -4710 5225
rect -6710 2740 -4710 2755
rect -4445 5225 -2445 5240
rect -4445 2755 -4430 5225
rect -2460 2755 -2445 5225
rect -4445 2740 -2445 2755
rect -2180 5225 -180 5240
rect -2180 2755 -2165 5225
rect -195 2755 -180 5225
rect -2180 2740 -180 2755
rect 85 5225 2085 5240
rect 85 2755 100 5225
rect 2070 2755 2085 5225
rect 85 2740 2085 2755
rect 2350 5225 4350 5240
rect 2350 2755 2365 5225
rect 4335 2755 4350 5225
rect 2350 2740 4350 2755
rect 4615 5225 6615 5240
rect 4615 2755 4630 5225
rect 6600 2755 6615 5225
rect 4615 2740 6615 2755
rect 6880 5225 8880 5240
rect 6880 2755 6895 5225
rect 8865 2755 8880 5225
rect 6880 2740 8880 2755
rect 9145 5225 11145 5240
rect 9145 2755 9160 5225
rect 11130 2755 11145 5225
rect 9145 2740 11145 2755
rect -11240 2565 -9240 2580
rect -11240 95 -11225 2565
rect -9255 95 -9240 2565
rect -11240 80 -9240 95
rect -8975 2565 -6975 2580
rect -8975 95 -8960 2565
rect -6990 95 -6975 2565
rect -8975 80 -6975 95
rect -6710 2565 -4710 2580
rect -6710 95 -6695 2565
rect -4725 95 -4710 2565
rect -6710 80 -4710 95
rect -4445 2565 -2445 2580
rect -4445 95 -4430 2565
rect -2460 95 -2445 2565
rect -4445 80 -2445 95
rect -2180 2565 -180 2580
rect -2180 95 -2165 2565
rect -195 95 -180 2565
rect -2180 80 -180 95
rect 85 2565 2085 2580
rect 85 95 100 2565
rect 2070 95 2085 2565
rect 85 80 2085 95
rect 2350 2565 4350 2580
rect 2350 95 2365 2565
rect 4335 95 4350 2565
rect 2350 80 4350 95
rect 4615 2565 6615 2580
rect 4615 95 4630 2565
rect 6600 95 6615 2565
rect 4615 80 6615 95
rect 6880 2565 8880 2580
rect 6880 95 6895 2565
rect 8865 95 8880 2565
rect 6880 80 8880 95
rect 9145 2565 11145 2580
rect 9145 95 9160 2565
rect 11130 95 11145 2565
rect 9145 80 11145 95
rect -11240 -95 -9240 -80
rect -11240 -2565 -11225 -95
rect -9255 -2565 -9240 -95
rect -11240 -2580 -9240 -2565
rect -8975 -95 -6975 -80
rect -8975 -2565 -8960 -95
rect -6990 -2565 -6975 -95
rect -8975 -2580 -6975 -2565
rect -6710 -95 -4710 -80
rect -6710 -2565 -6695 -95
rect -4725 -2565 -4710 -95
rect -6710 -2580 -4710 -2565
rect -4445 -95 -2445 -80
rect -4445 -2565 -4430 -95
rect -2460 -2565 -2445 -95
rect -4445 -2580 -2445 -2565
rect -2180 -95 -180 -80
rect -2180 -2565 -2165 -95
rect -195 -2565 -180 -95
rect -2180 -2580 -180 -2565
rect 85 -95 2085 -80
rect 85 -2565 100 -95
rect 2070 -2565 2085 -95
rect 85 -2580 2085 -2565
rect 2350 -95 4350 -80
rect 2350 -2565 2365 -95
rect 4335 -2565 4350 -95
rect 2350 -2580 4350 -2565
rect 4615 -95 6615 -80
rect 4615 -2565 4630 -95
rect 6600 -2565 6615 -95
rect 4615 -2580 6615 -2565
rect 6880 -95 8880 -80
rect 6880 -2565 6895 -95
rect 8865 -2565 8880 -95
rect 6880 -2580 8880 -2565
rect 9145 -95 11145 -80
rect 9145 -2565 9160 -95
rect 11130 -2565 11145 -95
rect 9145 -2580 11145 -2565
rect -11240 -2755 -9240 -2740
rect -11240 -5225 -11225 -2755
rect -9255 -5225 -9240 -2755
rect -11240 -5240 -9240 -5225
rect -8975 -2755 -6975 -2740
rect -8975 -5225 -8960 -2755
rect -6990 -5225 -6975 -2755
rect -8975 -5240 -6975 -5225
rect -6710 -2755 -4710 -2740
rect -6710 -5225 -6695 -2755
rect -4725 -5225 -4710 -2755
rect -6710 -5240 -4710 -5225
rect -4445 -2755 -2445 -2740
rect -4445 -5225 -4430 -2755
rect -2460 -5225 -2445 -2755
rect -4445 -5240 -2445 -5225
rect -2180 -2755 -180 -2740
rect -2180 -5225 -2165 -2755
rect -195 -5225 -180 -2755
rect -2180 -5240 -180 -5225
rect 85 -2755 2085 -2740
rect 85 -5225 100 -2755
rect 2070 -5225 2085 -2755
rect 85 -5240 2085 -5225
rect 2350 -2755 4350 -2740
rect 2350 -5225 2365 -2755
rect 4335 -5225 4350 -2755
rect 2350 -5240 4350 -5225
rect 4615 -2755 6615 -2740
rect 4615 -5225 4630 -2755
rect 6600 -5225 6615 -2755
rect 4615 -5240 6615 -5225
rect 6880 -2755 8880 -2740
rect 6880 -5225 6895 -2755
rect 8865 -5225 8880 -2755
rect 6880 -5240 8880 -5225
rect 9145 -2755 11145 -2740
rect 9145 -5225 9160 -2755
rect 11130 -5225 11145 -2755
rect 9145 -5240 11145 -5225
<< mimcapcontact >>
rect -11225 2755 -9255 5225
rect -8960 2755 -6990 5225
rect -6695 2755 -4725 5225
rect -4430 2755 -2460 5225
rect -2165 2755 -195 5225
rect 100 2755 2070 5225
rect 2365 2755 4335 5225
rect 4630 2755 6600 5225
rect 6895 2755 8865 5225
rect 9160 2755 11130 5225
rect -11225 95 -9255 2565
rect -8960 95 -6990 2565
rect -6695 95 -4725 2565
rect -4430 95 -2460 2565
rect -2165 95 -195 2565
rect 100 95 2070 2565
rect 2365 95 4335 2565
rect 4630 95 6600 2565
rect 6895 95 8865 2565
rect 9160 95 11130 2565
rect -11225 -2565 -9255 -95
rect -8960 -2565 -6990 -95
rect -6695 -2565 -4725 -95
rect -4430 -2565 -2460 -95
rect -2165 -2565 -195 -95
rect 100 -2565 2070 -95
rect 2365 -2565 4335 -95
rect 4630 -2565 6600 -95
rect 6895 -2565 8865 -95
rect 9160 -2565 11130 -95
rect -11225 -5225 -9255 -2755
rect -8960 -5225 -6990 -2755
rect -6695 -5225 -4725 -2755
rect -4430 -5225 -2460 -2755
rect -2165 -5225 -195 -2755
rect 100 -5225 2070 -2755
rect 2365 -5225 4335 -2755
rect 4630 -5225 6600 -2755
rect 6895 -5225 8865 -2755
rect 9160 -5225 11130 -2755
<< metal4 >>
rect -11290 5276 -9095 5290
rect -11290 5240 -9155 5276
rect -11290 2740 -11240 5240
rect -9240 2740 -9155 5240
rect -11290 2704 -9155 2740
rect -9105 2704 -9095 5276
rect -11290 2690 -9095 2704
rect -9025 5276 -6830 5290
rect -9025 5240 -6890 5276
rect -9025 2740 -8975 5240
rect -6975 2740 -6890 5240
rect -9025 2704 -6890 2740
rect -6840 2704 -6830 5276
rect -9025 2690 -6830 2704
rect -6760 5276 -4565 5290
rect -6760 5240 -4625 5276
rect -6760 2740 -6710 5240
rect -4710 2740 -4625 5240
rect -6760 2704 -4625 2740
rect -4575 2704 -4565 5276
rect -6760 2690 -4565 2704
rect -4495 5276 -2300 5290
rect -4495 5240 -2360 5276
rect -4495 2740 -4445 5240
rect -2445 2740 -2360 5240
rect -4495 2704 -2360 2740
rect -2310 2704 -2300 5276
rect -4495 2690 -2300 2704
rect -2230 5276 -35 5290
rect -2230 5240 -95 5276
rect -2230 2740 -2180 5240
rect -180 2740 -95 5240
rect -2230 2704 -95 2740
rect -45 2704 -35 5276
rect -2230 2690 -35 2704
rect 35 5276 2230 5290
rect 35 5240 2170 5276
rect 35 2740 85 5240
rect 2085 2740 2170 5240
rect 35 2704 2170 2740
rect 2220 2704 2230 5276
rect 35 2690 2230 2704
rect 2300 5276 4495 5290
rect 2300 5240 4435 5276
rect 2300 2740 2350 5240
rect 4350 2740 4435 5240
rect 2300 2704 4435 2740
rect 4485 2704 4495 5276
rect 2300 2690 4495 2704
rect 4565 5276 6760 5290
rect 4565 5240 6700 5276
rect 4565 2740 4615 5240
rect 6615 2740 6700 5240
rect 4565 2704 6700 2740
rect 6750 2704 6760 5276
rect 4565 2690 6760 2704
rect 6830 5276 9025 5290
rect 6830 5240 8965 5276
rect 6830 2740 6880 5240
rect 8880 2740 8965 5240
rect 6830 2704 8965 2740
rect 9015 2704 9025 5276
rect 6830 2690 9025 2704
rect 9095 5276 11290 5290
rect 9095 5240 11230 5276
rect 9095 2740 9145 5240
rect 11145 2740 11230 5240
rect 9095 2704 11230 2740
rect 11280 2704 11290 5276
rect 9095 2690 11290 2704
rect -11290 2616 -9095 2630
rect -11290 2580 -9155 2616
rect -11290 80 -11240 2580
rect -9240 80 -9155 2580
rect -11290 44 -9155 80
rect -9105 44 -9095 2616
rect -11290 30 -9095 44
rect -9025 2616 -6830 2630
rect -9025 2580 -6890 2616
rect -9025 80 -8975 2580
rect -6975 80 -6890 2580
rect -9025 44 -6890 80
rect -6840 44 -6830 2616
rect -9025 30 -6830 44
rect -6760 2616 -4565 2630
rect -6760 2580 -4625 2616
rect -6760 80 -6710 2580
rect -4710 80 -4625 2580
rect -6760 44 -4625 80
rect -4575 44 -4565 2616
rect -6760 30 -4565 44
rect -4495 2616 -2300 2630
rect -4495 2580 -2360 2616
rect -4495 80 -4445 2580
rect -2445 80 -2360 2580
rect -4495 44 -2360 80
rect -2310 44 -2300 2616
rect -4495 30 -2300 44
rect -2230 2616 -35 2630
rect -2230 2580 -95 2616
rect -2230 80 -2180 2580
rect -180 80 -95 2580
rect -2230 44 -95 80
rect -45 44 -35 2616
rect -2230 30 -35 44
rect 35 2616 2230 2630
rect 35 2580 2170 2616
rect 35 80 85 2580
rect 2085 80 2170 2580
rect 35 44 2170 80
rect 2220 44 2230 2616
rect 35 30 2230 44
rect 2300 2616 4495 2630
rect 2300 2580 4435 2616
rect 2300 80 2350 2580
rect 4350 80 4435 2580
rect 2300 44 4435 80
rect 4485 44 4495 2616
rect 2300 30 4495 44
rect 4565 2616 6760 2630
rect 4565 2580 6700 2616
rect 4565 80 4615 2580
rect 6615 80 6700 2580
rect 4565 44 6700 80
rect 6750 44 6760 2616
rect 4565 30 6760 44
rect 6830 2616 9025 2630
rect 6830 2580 8965 2616
rect 6830 80 6880 2580
rect 8880 80 8965 2580
rect 6830 44 8965 80
rect 9015 44 9025 2616
rect 6830 30 9025 44
rect 9095 2616 11290 2630
rect 9095 2580 11230 2616
rect 9095 80 9145 2580
rect 11145 80 11230 2580
rect 9095 44 11230 80
rect 11280 44 11290 2616
rect 9095 30 11290 44
rect -11290 -44 -9095 -30
rect -11290 -80 -9155 -44
rect -11290 -2580 -11240 -80
rect -9240 -2580 -9155 -80
rect -11290 -2616 -9155 -2580
rect -9105 -2616 -9095 -44
rect -11290 -2630 -9095 -2616
rect -9025 -44 -6830 -30
rect -9025 -80 -6890 -44
rect -9025 -2580 -8975 -80
rect -6975 -2580 -6890 -80
rect -9025 -2616 -6890 -2580
rect -6840 -2616 -6830 -44
rect -9025 -2630 -6830 -2616
rect -6760 -44 -4565 -30
rect -6760 -80 -4625 -44
rect -6760 -2580 -6710 -80
rect -4710 -2580 -4625 -80
rect -6760 -2616 -4625 -2580
rect -4575 -2616 -4565 -44
rect -6760 -2630 -4565 -2616
rect -4495 -44 -2300 -30
rect -4495 -80 -2360 -44
rect -4495 -2580 -4445 -80
rect -2445 -2580 -2360 -80
rect -4495 -2616 -2360 -2580
rect -2310 -2616 -2300 -44
rect -4495 -2630 -2300 -2616
rect -2230 -44 -35 -30
rect -2230 -80 -95 -44
rect -2230 -2580 -2180 -80
rect -180 -2580 -95 -80
rect -2230 -2616 -95 -2580
rect -45 -2616 -35 -44
rect -2230 -2630 -35 -2616
rect 35 -44 2230 -30
rect 35 -80 2170 -44
rect 35 -2580 85 -80
rect 2085 -2580 2170 -80
rect 35 -2616 2170 -2580
rect 2220 -2616 2230 -44
rect 35 -2630 2230 -2616
rect 2300 -44 4495 -30
rect 2300 -80 4435 -44
rect 2300 -2580 2350 -80
rect 4350 -2580 4435 -80
rect 2300 -2616 4435 -2580
rect 4485 -2616 4495 -44
rect 2300 -2630 4495 -2616
rect 4565 -44 6760 -30
rect 4565 -80 6700 -44
rect 4565 -2580 4615 -80
rect 6615 -2580 6700 -80
rect 4565 -2616 6700 -2580
rect 6750 -2616 6760 -44
rect 4565 -2630 6760 -2616
rect 6830 -44 9025 -30
rect 6830 -80 8965 -44
rect 6830 -2580 6880 -80
rect 8880 -2580 8965 -80
rect 6830 -2616 8965 -2580
rect 9015 -2616 9025 -44
rect 6830 -2630 9025 -2616
rect 9095 -44 11290 -30
rect 9095 -80 11230 -44
rect 9095 -2580 9145 -80
rect 11145 -2580 11230 -80
rect 9095 -2616 11230 -2580
rect 11280 -2616 11290 -44
rect 9095 -2630 11290 -2616
rect -11290 -2704 -9095 -2690
rect -11290 -2740 -9155 -2704
rect -11290 -5240 -11240 -2740
rect -9240 -5240 -9155 -2740
rect -11290 -5276 -9155 -5240
rect -9105 -5276 -9095 -2704
rect -11290 -5290 -9095 -5276
rect -9025 -2704 -6830 -2690
rect -9025 -2740 -6890 -2704
rect -9025 -5240 -8975 -2740
rect -6975 -5240 -6890 -2740
rect -9025 -5276 -6890 -5240
rect -6840 -5276 -6830 -2704
rect -9025 -5290 -6830 -5276
rect -6760 -2704 -4565 -2690
rect -6760 -2740 -4625 -2704
rect -6760 -5240 -6710 -2740
rect -4710 -5240 -4625 -2740
rect -6760 -5276 -4625 -5240
rect -4575 -5276 -4565 -2704
rect -6760 -5290 -4565 -5276
rect -4495 -2704 -2300 -2690
rect -4495 -2740 -2360 -2704
rect -4495 -5240 -4445 -2740
rect -2445 -5240 -2360 -2740
rect -4495 -5276 -2360 -5240
rect -2310 -5276 -2300 -2704
rect -4495 -5290 -2300 -5276
rect -2230 -2704 -35 -2690
rect -2230 -2740 -95 -2704
rect -2230 -5240 -2180 -2740
rect -180 -5240 -95 -2740
rect -2230 -5276 -95 -5240
rect -45 -5276 -35 -2704
rect -2230 -5290 -35 -5276
rect 35 -2704 2230 -2690
rect 35 -2740 2170 -2704
rect 35 -5240 85 -2740
rect 2085 -5240 2170 -2740
rect 35 -5276 2170 -5240
rect 2220 -5276 2230 -2704
rect 35 -5290 2230 -5276
rect 2300 -2704 4495 -2690
rect 2300 -2740 4435 -2704
rect 2300 -5240 2350 -2740
rect 4350 -5240 4435 -2740
rect 2300 -5276 4435 -5240
rect 4485 -5276 4495 -2704
rect 2300 -5290 4495 -5276
rect 4565 -2704 6760 -2690
rect 4565 -2740 6700 -2704
rect 4565 -5240 4615 -2740
rect 6615 -5240 6700 -2740
rect 4565 -5276 6700 -5240
rect 6750 -5276 6760 -2704
rect 4565 -5290 6760 -5276
rect 6830 -2704 9025 -2690
rect 6830 -2740 8965 -2704
rect 6830 -5240 6880 -2740
rect 8880 -5240 8965 -2740
rect 6830 -5276 8965 -5240
rect 9015 -5276 9025 -2704
rect 6830 -5290 9025 -5276
rect 9095 -2704 11290 -2690
rect 9095 -2740 11230 -2704
rect 9095 -5240 9145 -2740
rect 11145 -5240 11230 -2740
rect 9095 -5276 11230 -5240
rect 11280 -5276 11290 -2704
rect 9095 -5290 11290 -5276
<< viatp >>
rect -9155 2704 -9105 5276
rect -6890 2704 -6840 5276
rect -4625 2704 -4575 5276
rect -2360 2704 -2310 5276
rect -95 2704 -45 5276
rect 2170 2704 2220 5276
rect 4435 2704 4485 5276
rect 6700 2704 6750 5276
rect 8965 2704 9015 5276
rect 11230 2704 11280 5276
rect -9155 44 -9105 2616
rect -6890 44 -6840 2616
rect -4625 44 -4575 2616
rect -2360 44 -2310 2616
rect -95 44 -45 2616
rect 2170 44 2220 2616
rect 4435 44 4485 2616
rect 6700 44 6750 2616
rect 8965 44 9015 2616
rect 11230 44 11280 2616
rect -9155 -2616 -9105 -44
rect -6890 -2616 -6840 -44
rect -4625 -2616 -4575 -44
rect -2360 -2616 -2310 -44
rect -95 -2616 -45 -44
rect 2170 -2616 2220 -44
rect 4435 -2616 4485 -44
rect 6700 -2616 6750 -44
rect 8965 -2616 9015 -44
rect 11230 -2616 11280 -44
rect -9155 -5276 -9105 -2704
rect -6890 -5276 -6840 -2704
rect -4625 -5276 -4575 -2704
rect -2360 -5276 -2310 -2704
rect -95 -5276 -45 -2704
rect 2170 -5276 2220 -2704
rect 4435 -5276 4485 -2704
rect 6700 -5276 6750 -2704
rect 8965 -5276 9015 -2704
rect 11230 -5276 11280 -2704
<< metaltp >>
rect -10275 5225 -10205 5320
rect -9165 5276 -9095 5320
rect -10275 2565 -10205 2755
rect -9165 2704 -9155 5276
rect -9105 2704 -9095 5276
rect -8010 5225 -7940 5320
rect -6900 5276 -6830 5320
rect -9165 2616 -9095 2704
rect -10275 -95 -10205 95
rect -9165 44 -9155 2616
rect -9105 44 -9095 2616
rect -8010 2565 -7940 2755
rect -6900 2704 -6890 5276
rect -6840 2704 -6830 5276
rect -5745 5225 -5675 5320
rect -4635 5276 -4565 5320
rect -6900 2616 -6830 2704
rect -9165 -44 -9095 44
rect -10275 -2755 -10205 -2565
rect -9165 -2616 -9155 -44
rect -9105 -2616 -9095 -44
rect -8010 -95 -7940 95
rect -6900 44 -6890 2616
rect -6840 44 -6830 2616
rect -5745 2565 -5675 2755
rect -4635 2704 -4625 5276
rect -4575 2704 -4565 5276
rect -3480 5225 -3410 5320
rect -2370 5276 -2300 5320
rect -4635 2616 -4565 2704
rect -6900 -44 -6830 44
rect -9165 -2704 -9095 -2616
rect -10275 -5320 -10205 -5225
rect -9165 -5276 -9155 -2704
rect -9105 -5276 -9095 -2704
rect -8010 -2755 -7940 -2565
rect -6900 -2616 -6890 -44
rect -6840 -2616 -6830 -44
rect -5745 -95 -5675 95
rect -4635 44 -4625 2616
rect -4575 44 -4565 2616
rect -3480 2565 -3410 2755
rect -2370 2704 -2360 5276
rect -2310 2704 -2300 5276
rect -1215 5225 -1145 5320
rect -105 5276 -35 5320
rect -2370 2616 -2300 2704
rect -4635 -44 -4565 44
rect -6900 -2704 -6830 -2616
rect -9165 -5320 -9095 -5276
rect -8010 -5320 -7940 -5225
rect -6900 -5276 -6890 -2704
rect -6840 -5276 -6830 -2704
rect -5745 -2755 -5675 -2565
rect -4635 -2616 -4625 -44
rect -4575 -2616 -4565 -44
rect -3480 -95 -3410 95
rect -2370 44 -2360 2616
rect -2310 44 -2300 2616
rect -1215 2565 -1145 2755
rect -105 2704 -95 5276
rect -45 2704 -35 5276
rect 1050 5225 1120 5320
rect 2160 5276 2230 5320
rect -105 2616 -35 2704
rect -2370 -44 -2300 44
rect -4635 -2704 -4565 -2616
rect -6900 -5320 -6830 -5276
rect -5745 -5320 -5675 -5225
rect -4635 -5276 -4625 -2704
rect -4575 -5276 -4565 -2704
rect -3480 -2755 -3410 -2565
rect -2370 -2616 -2360 -44
rect -2310 -2616 -2300 -44
rect -1215 -95 -1145 95
rect -105 44 -95 2616
rect -45 44 -35 2616
rect 1050 2565 1120 2755
rect 2160 2704 2170 5276
rect 2220 2704 2230 5276
rect 3315 5225 3385 5320
rect 4425 5276 4495 5320
rect 2160 2616 2230 2704
rect -105 -44 -35 44
rect -2370 -2704 -2300 -2616
rect -4635 -5320 -4565 -5276
rect -3480 -5320 -3410 -5225
rect -2370 -5276 -2360 -2704
rect -2310 -5276 -2300 -2704
rect -1215 -2755 -1145 -2565
rect -105 -2616 -95 -44
rect -45 -2616 -35 -44
rect 1050 -95 1120 95
rect 2160 44 2170 2616
rect 2220 44 2230 2616
rect 3315 2565 3385 2755
rect 4425 2704 4435 5276
rect 4485 2704 4495 5276
rect 5580 5225 5650 5320
rect 6690 5276 6760 5320
rect 4425 2616 4495 2704
rect 2160 -44 2230 44
rect -105 -2704 -35 -2616
rect -2370 -5320 -2300 -5276
rect -1215 -5320 -1145 -5225
rect -105 -5276 -95 -2704
rect -45 -5276 -35 -2704
rect 1050 -2755 1120 -2565
rect 2160 -2616 2170 -44
rect 2220 -2616 2230 -44
rect 3315 -95 3385 95
rect 4425 44 4435 2616
rect 4485 44 4495 2616
rect 5580 2565 5650 2755
rect 6690 2704 6700 5276
rect 6750 2704 6760 5276
rect 7845 5225 7915 5320
rect 8955 5276 9025 5320
rect 6690 2616 6760 2704
rect 4425 -44 4495 44
rect 2160 -2704 2230 -2616
rect -105 -5320 -35 -5276
rect 1050 -5320 1120 -5225
rect 2160 -5276 2170 -2704
rect 2220 -5276 2230 -2704
rect 3315 -2755 3385 -2565
rect 4425 -2616 4435 -44
rect 4485 -2616 4495 -44
rect 5580 -95 5650 95
rect 6690 44 6700 2616
rect 6750 44 6760 2616
rect 7845 2565 7915 2755
rect 8955 2704 8965 5276
rect 9015 2704 9025 5276
rect 10110 5225 10180 5320
rect 11220 5276 11290 5320
rect 8955 2616 9025 2704
rect 6690 -44 6760 44
rect 4425 -2704 4495 -2616
rect 2160 -5320 2230 -5276
rect 3315 -5320 3385 -5225
rect 4425 -5276 4435 -2704
rect 4485 -5276 4495 -2704
rect 5580 -2755 5650 -2565
rect 6690 -2616 6700 -44
rect 6750 -2616 6760 -44
rect 7845 -95 7915 95
rect 8955 44 8965 2616
rect 9015 44 9025 2616
rect 10110 2565 10180 2755
rect 11220 2704 11230 5276
rect 11280 2704 11290 5276
rect 11220 2616 11290 2704
rect 8955 -44 9025 44
rect 6690 -2704 6760 -2616
rect 4425 -5320 4495 -5276
rect 5580 -5320 5650 -5225
rect 6690 -5276 6700 -2704
rect 6750 -5276 6760 -2704
rect 7845 -2755 7915 -2565
rect 8955 -2616 8965 -44
rect 9015 -2616 9025 -44
rect 10110 -95 10180 95
rect 11220 44 11230 2616
rect 11280 44 11290 2616
rect 11220 -44 11290 44
rect 8955 -2704 9025 -2616
rect 6690 -5320 6760 -5276
rect 7845 -5320 7915 -5225
rect 8955 -5276 8965 -2704
rect 9015 -5276 9025 -2704
rect 10110 -2755 10180 -2565
rect 11220 -2616 11230 -44
rect 11280 -2616 11290 -44
rect 11220 -2704 11290 -2616
rect 8955 -5320 9025 -5276
rect 10110 -5320 10180 -5225
rect 11220 -5276 11230 -2704
rect 11280 -5276 11290 -2704
rect 11220 -5320 11290 -5276
<< boundary >>
rect -11290 2690 -9190 5290
rect -9025 2690 -6925 5290
rect -6760 2690 -4660 5290
rect -4495 2690 -2395 5290
rect -2230 2690 -130 5290
rect 35 2690 2135 5290
rect 2300 2690 4400 5290
rect 4565 2690 6665 5290
rect 6830 2690 8930 5290
rect 9095 2690 11195 5290
rect -11290 30 -9190 2630
rect -9025 30 -6925 2630
rect -6760 30 -4660 2630
rect -4495 30 -2395 2630
rect -2230 30 -130 2630
rect 35 30 2135 2630
rect 2300 30 4400 2630
rect 4565 30 6665 2630
rect 6830 30 8930 2630
rect 9095 30 11195 2630
rect -11290 -2630 -9190 -30
rect -9025 -2630 -6925 -30
rect -6760 -2630 -4660 -30
rect -4495 -2630 -2395 -30
rect -2230 -2630 -130 -30
rect 35 -2630 2135 -30
rect 2300 -2630 4400 -30
rect 4565 -2630 6665 -30
rect 6830 -2630 8930 -30
rect 9095 -2630 11195 -30
rect -11290 -5290 -9190 -2690
rect -9025 -5290 -6925 -2690
rect -6760 -5290 -4660 -2690
rect -4495 -5290 -2395 -2690
rect -2230 -5290 -130 -2690
rect 35 -5290 2135 -2690
rect 2300 -5290 4400 -2690
rect 4565 -5290 6665 -2690
rect 6830 -5290 8930 -2690
rect 9095 -5290 11195 -2690
<< properties >>
string parameters w 20.00 l 25.00 val 515.299 carea 1.00 cperi 0.17 nx 10 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
