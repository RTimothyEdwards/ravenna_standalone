magic
tech EFXH018D
timestamp 1533305873
<< mimcap >>
rect -4445 7465 -2445 7480
rect -4445 5495 -4430 7465
rect -2460 5495 -2445 7465
rect -4445 5480 -2445 5495
rect -2180 7465 -180 7480
rect -2180 5495 -2165 7465
rect -195 5495 -180 7465
rect -2180 5480 -180 5495
rect 85 7465 2085 7480
rect 85 5495 100 7465
rect 2070 5495 2085 7465
rect 85 5480 2085 5495
rect 2350 7465 4350 7480
rect 2350 5495 2365 7465
rect 4335 5495 4350 7465
rect 2350 5480 4350 5495
rect -4445 5305 -2445 5320
rect -4445 3335 -4430 5305
rect -2460 3335 -2445 5305
rect -4445 3320 -2445 3335
rect -2180 5305 -180 5320
rect -2180 3335 -2165 5305
rect -195 3335 -180 5305
rect -2180 3320 -180 3335
rect 85 5305 2085 5320
rect 85 3335 100 5305
rect 2070 3335 2085 5305
rect 85 3320 2085 3335
rect 2350 5305 4350 5320
rect 2350 3335 2365 5305
rect 4335 3335 4350 5305
rect 2350 3320 4350 3335
rect -4445 3145 -2445 3160
rect -4445 1175 -4430 3145
rect -2460 1175 -2445 3145
rect -4445 1160 -2445 1175
rect -2180 3145 -180 3160
rect -2180 1175 -2165 3145
rect -195 1175 -180 3145
rect -2180 1160 -180 1175
rect 85 3145 2085 3160
rect 85 1175 100 3145
rect 2070 1175 2085 3145
rect 85 1160 2085 1175
rect 2350 3145 4350 3160
rect 2350 1175 2365 3145
rect 4335 1175 4350 3145
rect 2350 1160 4350 1175
rect -4445 985 -2445 1000
rect -4445 -985 -4430 985
rect -2460 -985 -2445 985
rect -4445 -1000 -2445 -985
rect -2180 985 -180 1000
rect -2180 -985 -2165 985
rect -195 -985 -180 985
rect -2180 -1000 -180 -985
rect 85 985 2085 1000
rect 85 -985 100 985
rect 2070 -985 2085 985
rect 85 -1000 2085 -985
rect 2350 985 4350 1000
rect 2350 -985 2365 985
rect 4335 -985 4350 985
rect 2350 -1000 4350 -985
rect -4445 -1175 -2445 -1160
rect -4445 -3145 -4430 -1175
rect -2460 -3145 -2445 -1175
rect -4445 -3160 -2445 -3145
rect -2180 -1175 -180 -1160
rect -2180 -3145 -2165 -1175
rect -195 -3145 -180 -1175
rect -2180 -3160 -180 -3145
rect 85 -1175 2085 -1160
rect 85 -3145 100 -1175
rect 2070 -3145 2085 -1175
rect 85 -3160 2085 -3145
rect 2350 -1175 4350 -1160
rect 2350 -3145 2365 -1175
rect 4335 -3145 4350 -1175
rect 2350 -3160 4350 -3145
rect -4445 -3335 -2445 -3320
rect -4445 -5305 -4430 -3335
rect -2460 -5305 -2445 -3335
rect -4445 -5320 -2445 -5305
rect -2180 -3335 -180 -3320
rect -2180 -5305 -2165 -3335
rect -195 -5305 -180 -3335
rect -2180 -5320 -180 -5305
rect 85 -3335 2085 -3320
rect 85 -5305 100 -3335
rect 2070 -5305 2085 -3335
rect 85 -5320 2085 -5305
rect 2350 -3335 4350 -3320
rect 2350 -5305 2365 -3335
rect 4335 -5305 4350 -3335
rect 2350 -5320 4350 -5305
rect -4445 -5495 -2445 -5480
rect -4445 -7465 -4430 -5495
rect -2460 -7465 -2445 -5495
rect -4445 -7480 -2445 -7465
rect -2180 -5495 -180 -5480
rect -2180 -7465 -2165 -5495
rect -195 -7465 -180 -5495
rect -2180 -7480 -180 -7465
rect 85 -5495 2085 -5480
rect 85 -7465 100 -5495
rect 2070 -7465 2085 -5495
rect 85 -7480 2085 -7465
rect 2350 -5495 4350 -5480
rect 2350 -7465 2365 -5495
rect 4335 -7465 4350 -5495
rect 2350 -7480 4350 -7465
<< mimcapcontact >>
rect -4430 5495 -2460 7465
rect -2165 5495 -195 7465
rect 100 5495 2070 7465
rect 2365 5495 4335 7465
rect -4430 3335 -2460 5305
rect -2165 3335 -195 5305
rect 100 3335 2070 5305
rect 2365 3335 4335 5305
rect -4430 1175 -2460 3145
rect -2165 1175 -195 3145
rect 100 1175 2070 3145
rect 2365 1175 4335 3145
rect -4430 -985 -2460 985
rect -2165 -985 -195 985
rect 100 -985 2070 985
rect 2365 -985 4335 985
rect -4430 -3145 -2460 -1175
rect -2165 -3145 -195 -1175
rect 100 -3145 2070 -1175
rect 2365 -3145 4335 -1175
rect -4430 -5305 -2460 -3335
rect -2165 -5305 -195 -3335
rect 100 -5305 2070 -3335
rect 2365 -5305 4335 -3335
rect -4430 -7465 -2460 -5495
rect -2165 -7465 -195 -5495
rect 100 -7465 2070 -5495
rect 2365 -7465 4335 -5495
<< metal4 >>
rect -4495 7516 -2300 7530
rect -4495 7480 -2360 7516
rect -4495 5480 -4445 7480
rect -2445 5480 -2360 7480
rect -4495 5444 -2360 5480
rect -2310 5444 -2300 7516
rect -4495 5430 -2300 5444
rect -2230 7516 -35 7530
rect -2230 7480 -95 7516
rect -2230 5480 -2180 7480
rect -180 5480 -95 7480
rect -2230 5444 -95 5480
rect -45 5444 -35 7516
rect -2230 5430 -35 5444
rect 35 7516 2230 7530
rect 35 7480 2170 7516
rect 35 5480 85 7480
rect 2085 5480 2170 7480
rect 35 5444 2170 5480
rect 2220 5444 2230 7516
rect 35 5430 2230 5444
rect 2300 7516 4495 7530
rect 2300 7480 4435 7516
rect 2300 5480 2350 7480
rect 4350 5480 4435 7480
rect 2300 5444 4435 5480
rect 4485 5444 4495 7516
rect 2300 5430 4495 5444
rect -4495 5356 -2300 5370
rect -4495 5320 -2360 5356
rect -4495 3320 -4445 5320
rect -2445 3320 -2360 5320
rect -4495 3284 -2360 3320
rect -2310 3284 -2300 5356
rect -4495 3270 -2300 3284
rect -2230 5356 -35 5370
rect -2230 5320 -95 5356
rect -2230 3320 -2180 5320
rect -180 3320 -95 5320
rect -2230 3284 -95 3320
rect -45 3284 -35 5356
rect -2230 3270 -35 3284
rect 35 5356 2230 5370
rect 35 5320 2170 5356
rect 35 3320 85 5320
rect 2085 3320 2170 5320
rect 35 3284 2170 3320
rect 2220 3284 2230 5356
rect 35 3270 2230 3284
rect 2300 5356 4495 5370
rect 2300 5320 4435 5356
rect 2300 3320 2350 5320
rect 4350 3320 4435 5320
rect 2300 3284 4435 3320
rect 4485 3284 4495 5356
rect 2300 3270 4495 3284
rect -4495 3196 -2300 3210
rect -4495 3160 -2360 3196
rect -4495 1160 -4445 3160
rect -2445 1160 -2360 3160
rect -4495 1124 -2360 1160
rect -2310 1124 -2300 3196
rect -4495 1110 -2300 1124
rect -2230 3196 -35 3210
rect -2230 3160 -95 3196
rect -2230 1160 -2180 3160
rect -180 1160 -95 3160
rect -2230 1124 -95 1160
rect -45 1124 -35 3196
rect -2230 1110 -35 1124
rect 35 3196 2230 3210
rect 35 3160 2170 3196
rect 35 1160 85 3160
rect 2085 1160 2170 3160
rect 35 1124 2170 1160
rect 2220 1124 2230 3196
rect 35 1110 2230 1124
rect 2300 3196 4495 3210
rect 2300 3160 4435 3196
rect 2300 1160 2350 3160
rect 4350 1160 4435 3160
rect 2300 1124 4435 1160
rect 4485 1124 4495 3196
rect 2300 1110 4495 1124
rect -4495 1036 -2300 1050
rect -4495 1000 -2360 1036
rect -4495 -1000 -4445 1000
rect -2445 -1000 -2360 1000
rect -4495 -1036 -2360 -1000
rect -2310 -1036 -2300 1036
rect -4495 -1050 -2300 -1036
rect -2230 1036 -35 1050
rect -2230 1000 -95 1036
rect -2230 -1000 -2180 1000
rect -180 -1000 -95 1000
rect -2230 -1036 -95 -1000
rect -45 -1036 -35 1036
rect -2230 -1050 -35 -1036
rect 35 1036 2230 1050
rect 35 1000 2170 1036
rect 35 -1000 85 1000
rect 2085 -1000 2170 1000
rect 35 -1036 2170 -1000
rect 2220 -1036 2230 1036
rect 35 -1050 2230 -1036
rect 2300 1036 4495 1050
rect 2300 1000 4435 1036
rect 2300 -1000 2350 1000
rect 4350 -1000 4435 1000
rect 2300 -1036 4435 -1000
rect 4485 -1036 4495 1036
rect 2300 -1050 4495 -1036
rect -4495 -1124 -2300 -1110
rect -4495 -1160 -2360 -1124
rect -4495 -3160 -4445 -1160
rect -2445 -3160 -2360 -1160
rect -4495 -3196 -2360 -3160
rect -2310 -3196 -2300 -1124
rect -4495 -3210 -2300 -3196
rect -2230 -1124 -35 -1110
rect -2230 -1160 -95 -1124
rect -2230 -3160 -2180 -1160
rect -180 -3160 -95 -1160
rect -2230 -3196 -95 -3160
rect -45 -3196 -35 -1124
rect -2230 -3210 -35 -3196
rect 35 -1124 2230 -1110
rect 35 -1160 2170 -1124
rect 35 -3160 85 -1160
rect 2085 -3160 2170 -1160
rect 35 -3196 2170 -3160
rect 2220 -3196 2230 -1124
rect 35 -3210 2230 -3196
rect 2300 -1124 4495 -1110
rect 2300 -1160 4435 -1124
rect 2300 -3160 2350 -1160
rect 4350 -3160 4435 -1160
rect 2300 -3196 4435 -3160
rect 4485 -3196 4495 -1124
rect 2300 -3210 4495 -3196
rect -4495 -3284 -2300 -3270
rect -4495 -3320 -2360 -3284
rect -4495 -5320 -4445 -3320
rect -2445 -5320 -2360 -3320
rect -4495 -5356 -2360 -5320
rect -2310 -5356 -2300 -3284
rect -4495 -5370 -2300 -5356
rect -2230 -3284 -35 -3270
rect -2230 -3320 -95 -3284
rect -2230 -5320 -2180 -3320
rect -180 -5320 -95 -3320
rect -2230 -5356 -95 -5320
rect -45 -5356 -35 -3284
rect -2230 -5370 -35 -5356
rect 35 -3284 2230 -3270
rect 35 -3320 2170 -3284
rect 35 -5320 85 -3320
rect 2085 -5320 2170 -3320
rect 35 -5356 2170 -5320
rect 2220 -5356 2230 -3284
rect 35 -5370 2230 -5356
rect 2300 -3284 4495 -3270
rect 2300 -3320 4435 -3284
rect 2300 -5320 2350 -3320
rect 4350 -5320 4435 -3320
rect 2300 -5356 4435 -5320
rect 4485 -5356 4495 -3284
rect 2300 -5370 4495 -5356
rect -4495 -5444 -2300 -5430
rect -4495 -5480 -2360 -5444
rect -4495 -7480 -4445 -5480
rect -2445 -7480 -2360 -5480
rect -4495 -7516 -2360 -7480
rect -2310 -7516 -2300 -5444
rect -4495 -7530 -2300 -7516
rect -2230 -5444 -35 -5430
rect -2230 -5480 -95 -5444
rect -2230 -7480 -2180 -5480
rect -180 -7480 -95 -5480
rect -2230 -7516 -95 -7480
rect -45 -7516 -35 -5444
rect -2230 -7530 -35 -7516
rect 35 -5444 2230 -5430
rect 35 -5480 2170 -5444
rect 35 -7480 85 -5480
rect 2085 -7480 2170 -5480
rect 35 -7516 2170 -7480
rect 2220 -7516 2230 -5444
rect 35 -7530 2230 -7516
rect 2300 -5444 4495 -5430
rect 2300 -5480 4435 -5444
rect 2300 -7480 2350 -5480
rect 4350 -7480 4435 -5480
rect 2300 -7516 4435 -7480
rect 4485 -7516 4495 -5444
rect 2300 -7530 4495 -7516
<< viatp >>
rect -2360 5444 -2310 7516
rect -95 5444 -45 7516
rect 2170 5444 2220 7516
rect 4435 5444 4485 7516
rect -2360 3284 -2310 5356
rect -95 3284 -45 5356
rect 2170 3284 2220 5356
rect 4435 3284 4485 5356
rect -2360 1124 -2310 3196
rect -95 1124 -45 3196
rect 2170 1124 2220 3196
rect 4435 1124 4485 3196
rect -2360 -1036 -2310 1036
rect -95 -1036 -45 1036
rect 2170 -1036 2220 1036
rect 4435 -1036 4485 1036
rect -2360 -3196 -2310 -1124
rect -95 -3196 -45 -1124
rect 2170 -3196 2220 -1124
rect 4435 -3196 4485 -1124
rect -2360 -5356 -2310 -3284
rect -95 -5356 -45 -3284
rect 2170 -5356 2220 -3284
rect 4435 -5356 4485 -3284
rect -2360 -7516 -2310 -5444
rect -95 -7516 -45 -5444
rect 2170 -7516 2220 -5444
rect 4435 -7516 4485 -5444
<< metaltp >>
rect -3480 7465 -3410 7560
rect -2370 7516 -2300 7560
rect -3480 5305 -3410 5495
rect -2370 5444 -2360 7516
rect -2310 5444 -2300 7516
rect -1215 7465 -1145 7560
rect -105 7516 -35 7560
rect -2370 5356 -2300 5444
rect -3480 3145 -3410 3335
rect -2370 3284 -2360 5356
rect -2310 3284 -2300 5356
rect -1215 5305 -1145 5495
rect -105 5444 -95 7516
rect -45 5444 -35 7516
rect 1050 7465 1120 7560
rect 2160 7516 2230 7560
rect -105 5356 -35 5444
rect -2370 3196 -2300 3284
rect -3480 985 -3410 1175
rect -2370 1124 -2360 3196
rect -2310 1124 -2300 3196
rect -1215 3145 -1145 3335
rect -105 3284 -95 5356
rect -45 3284 -35 5356
rect 1050 5305 1120 5495
rect 2160 5444 2170 7516
rect 2220 5444 2230 7516
rect 3315 7465 3385 7560
rect 4425 7516 4495 7560
rect 2160 5356 2230 5444
rect -105 3196 -35 3284
rect -2370 1036 -2300 1124
rect -3480 -1175 -3410 -985
rect -2370 -1036 -2360 1036
rect -2310 -1036 -2300 1036
rect -1215 985 -1145 1175
rect -105 1124 -95 3196
rect -45 1124 -35 3196
rect 1050 3145 1120 3335
rect 2160 3284 2170 5356
rect 2220 3284 2230 5356
rect 3315 5305 3385 5495
rect 4425 5444 4435 7516
rect 4485 5444 4495 7516
rect 4425 5356 4495 5444
rect 2160 3196 2230 3284
rect -105 1036 -35 1124
rect -2370 -1124 -2300 -1036
rect -3480 -3335 -3410 -3145
rect -2370 -3196 -2360 -1124
rect -2310 -3196 -2300 -1124
rect -1215 -1175 -1145 -985
rect -105 -1036 -95 1036
rect -45 -1036 -35 1036
rect 1050 985 1120 1175
rect 2160 1124 2170 3196
rect 2220 1124 2230 3196
rect 3315 3145 3385 3335
rect 4425 3284 4435 5356
rect 4485 3284 4495 5356
rect 4425 3196 4495 3284
rect 2160 1036 2230 1124
rect -105 -1124 -35 -1036
rect -2370 -3284 -2300 -3196
rect -3480 -5495 -3410 -5305
rect -2370 -5356 -2360 -3284
rect -2310 -5356 -2300 -3284
rect -1215 -3335 -1145 -3145
rect -105 -3196 -95 -1124
rect -45 -3196 -35 -1124
rect 1050 -1175 1120 -985
rect 2160 -1036 2170 1036
rect 2220 -1036 2230 1036
rect 3315 985 3385 1175
rect 4425 1124 4435 3196
rect 4485 1124 4495 3196
rect 4425 1036 4495 1124
rect 2160 -1124 2230 -1036
rect -105 -3284 -35 -3196
rect -2370 -5444 -2300 -5356
rect -3480 -7560 -3410 -7465
rect -2370 -7516 -2360 -5444
rect -2310 -7516 -2300 -5444
rect -1215 -5495 -1145 -5305
rect -105 -5356 -95 -3284
rect -45 -5356 -35 -3284
rect 1050 -3335 1120 -3145
rect 2160 -3196 2170 -1124
rect 2220 -3196 2230 -1124
rect 3315 -1175 3385 -985
rect 4425 -1036 4435 1036
rect 4485 -1036 4495 1036
rect 4425 -1124 4495 -1036
rect 2160 -3284 2230 -3196
rect -105 -5444 -35 -5356
rect -2370 -7560 -2300 -7516
rect -1215 -7560 -1145 -7465
rect -105 -7516 -95 -5444
rect -45 -7516 -35 -5444
rect 1050 -5495 1120 -5305
rect 2160 -5356 2170 -3284
rect 2220 -5356 2230 -3284
rect 3315 -3335 3385 -3145
rect 4425 -3196 4435 -1124
rect 4485 -3196 4495 -1124
rect 4425 -3284 4495 -3196
rect 2160 -5444 2230 -5356
rect -105 -7560 -35 -7516
rect 1050 -7560 1120 -7465
rect 2160 -7516 2170 -5444
rect 2220 -7516 2230 -5444
rect 3315 -5495 3385 -5305
rect 4425 -5356 4435 -3284
rect 4485 -5356 4495 -3284
rect 4425 -5444 4495 -5356
rect 2160 -7560 2230 -7516
rect 3315 -7560 3385 -7465
rect 4425 -7516 4435 -5444
rect 4485 -7516 4495 -5444
rect 4425 -7560 4495 -7516
<< boundary >>
rect -4495 5430 -2395 7530
rect -2230 5430 -130 7530
rect 35 5430 2135 7530
rect 2300 5430 4400 7530
rect -4495 3270 -2395 5370
rect -2230 3270 -130 5370
rect 35 3270 2135 5370
rect 2300 3270 4400 5370
rect -4495 1110 -2395 3210
rect -2230 1110 -130 3210
rect 35 1110 2135 3210
rect 2300 1110 4400 3210
rect -4495 -1050 -2395 1050
rect -2230 -1050 -130 1050
rect 35 -1050 2135 1050
rect 2300 -1050 4400 1050
rect -4495 -3210 -2395 -1110
rect -2230 -3210 -130 -1110
rect 35 -3210 2135 -1110
rect 2300 -3210 4400 -1110
rect -4495 -5370 -2395 -3270
rect -2230 -5370 -130 -3270
rect 35 -5370 2135 -3270
rect 2300 -5370 4400 -3270
rect -4495 -7530 -2395 -5430
rect -2230 -7530 -130 -5430
rect 35 -7530 2135 -5430
rect 2300 -7530 4400 -5430
<< properties >>
string parameters w 20.00 l 20.00 val 413.6 carea 1.00 cperi 0.17 nx 4 ny 7 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
