magic
tech EFXH018D
timestamp 1565723183
<< mimcap >>
rect -13505 7465 -11505 7480
rect -13505 5495 -13490 7465
rect -11520 5495 -11505 7465
rect -13505 5480 -11505 5495
rect -11240 7465 -9240 7480
rect -11240 5495 -11225 7465
rect -9255 5495 -9240 7465
rect -11240 5480 -9240 5495
rect -8975 7465 -6975 7480
rect -8975 5495 -8960 7465
rect -6990 5495 -6975 7465
rect -8975 5480 -6975 5495
rect -6710 7465 -4710 7480
rect -6710 5495 -6695 7465
rect -4725 5495 -4710 7465
rect -6710 5480 -4710 5495
rect -4445 7465 -2445 7480
rect -4445 5495 -4430 7465
rect -2460 5495 -2445 7465
rect -4445 5480 -2445 5495
rect -2180 7465 -180 7480
rect -2180 5495 -2165 7465
rect -195 5495 -180 7465
rect -2180 5480 -180 5495
rect 85 7465 2085 7480
rect 85 5495 100 7465
rect 2070 5495 2085 7465
rect 85 5480 2085 5495
rect 2350 7465 4350 7480
rect 2350 5495 2365 7465
rect 4335 5495 4350 7465
rect 2350 5480 4350 5495
rect 4615 7465 6615 7480
rect 4615 5495 4630 7465
rect 6600 5495 6615 7465
rect 4615 5480 6615 5495
rect 6880 7465 8880 7480
rect 6880 5495 6895 7465
rect 8865 5495 8880 7465
rect 6880 5480 8880 5495
rect 9145 7465 11145 7480
rect 9145 5495 9160 7465
rect 11130 5495 11145 7465
rect 9145 5480 11145 5495
rect 11410 7465 13410 7480
rect 11410 5495 11425 7465
rect 13395 5495 13410 7465
rect 11410 5480 13410 5495
rect -13505 5305 -11505 5320
rect -13505 3335 -13490 5305
rect -11520 3335 -11505 5305
rect -13505 3320 -11505 3335
rect -11240 5305 -9240 5320
rect -11240 3335 -11225 5305
rect -9255 3335 -9240 5305
rect -11240 3320 -9240 3335
rect -8975 5305 -6975 5320
rect -8975 3335 -8960 5305
rect -6990 3335 -6975 5305
rect -8975 3320 -6975 3335
rect -6710 5305 -4710 5320
rect -6710 3335 -6695 5305
rect -4725 3335 -4710 5305
rect -6710 3320 -4710 3335
rect -4445 5305 -2445 5320
rect -4445 3335 -4430 5305
rect -2460 3335 -2445 5305
rect -4445 3320 -2445 3335
rect -2180 5305 -180 5320
rect -2180 3335 -2165 5305
rect -195 3335 -180 5305
rect -2180 3320 -180 3335
rect 85 5305 2085 5320
rect 85 3335 100 5305
rect 2070 3335 2085 5305
rect 85 3320 2085 3335
rect 2350 5305 4350 5320
rect 2350 3335 2365 5305
rect 4335 3335 4350 5305
rect 2350 3320 4350 3335
rect 4615 5305 6615 5320
rect 4615 3335 4630 5305
rect 6600 3335 6615 5305
rect 4615 3320 6615 3335
rect 6880 5305 8880 5320
rect 6880 3335 6895 5305
rect 8865 3335 8880 5305
rect 6880 3320 8880 3335
rect 9145 5305 11145 5320
rect 9145 3335 9160 5305
rect 11130 3335 11145 5305
rect 9145 3320 11145 3335
rect 11410 5305 13410 5320
rect 11410 3335 11425 5305
rect 13395 3335 13410 5305
rect 11410 3320 13410 3335
rect -13505 3145 -11505 3160
rect -13505 1175 -13490 3145
rect -11520 1175 -11505 3145
rect -13505 1160 -11505 1175
rect -11240 3145 -9240 3160
rect -11240 1175 -11225 3145
rect -9255 1175 -9240 3145
rect -11240 1160 -9240 1175
rect -8975 3145 -6975 3160
rect -8975 1175 -8960 3145
rect -6990 1175 -6975 3145
rect -8975 1160 -6975 1175
rect -6710 3145 -4710 3160
rect -6710 1175 -6695 3145
rect -4725 1175 -4710 3145
rect -6710 1160 -4710 1175
rect -4445 3145 -2445 3160
rect -4445 1175 -4430 3145
rect -2460 1175 -2445 3145
rect -4445 1160 -2445 1175
rect -2180 3145 -180 3160
rect -2180 1175 -2165 3145
rect -195 1175 -180 3145
rect -2180 1160 -180 1175
rect 85 3145 2085 3160
rect 85 1175 100 3145
rect 2070 1175 2085 3145
rect 85 1160 2085 1175
rect 2350 3145 4350 3160
rect 2350 1175 2365 3145
rect 4335 1175 4350 3145
rect 2350 1160 4350 1175
rect 4615 3145 6615 3160
rect 4615 1175 4630 3145
rect 6600 1175 6615 3145
rect 4615 1160 6615 1175
rect 6880 3145 8880 3160
rect 6880 1175 6895 3145
rect 8865 1175 8880 3145
rect 6880 1160 8880 1175
rect 9145 3145 11145 3160
rect 9145 1175 9160 3145
rect 11130 1175 11145 3145
rect 9145 1160 11145 1175
rect 11410 3145 13410 3160
rect 11410 1175 11425 3145
rect 13395 1175 13410 3145
rect 11410 1160 13410 1175
rect -13505 985 -11505 1000
rect -13505 -985 -13490 985
rect -11520 -985 -11505 985
rect -13505 -1000 -11505 -985
rect -11240 985 -9240 1000
rect -11240 -985 -11225 985
rect -9255 -985 -9240 985
rect -11240 -1000 -9240 -985
rect -8975 985 -6975 1000
rect -8975 -985 -8960 985
rect -6990 -985 -6975 985
rect -8975 -1000 -6975 -985
rect -6710 985 -4710 1000
rect -6710 -985 -6695 985
rect -4725 -985 -4710 985
rect -6710 -1000 -4710 -985
rect -4445 985 -2445 1000
rect -4445 -985 -4430 985
rect -2460 -985 -2445 985
rect -4445 -1000 -2445 -985
rect -2180 985 -180 1000
rect -2180 -985 -2165 985
rect -195 -985 -180 985
rect -2180 -1000 -180 -985
rect 85 985 2085 1000
rect 85 -985 100 985
rect 2070 -985 2085 985
rect 85 -1000 2085 -985
rect 2350 985 4350 1000
rect 2350 -985 2365 985
rect 4335 -985 4350 985
rect 2350 -1000 4350 -985
rect 4615 985 6615 1000
rect 4615 -985 4630 985
rect 6600 -985 6615 985
rect 4615 -1000 6615 -985
rect 6880 985 8880 1000
rect 6880 -985 6895 985
rect 8865 -985 8880 985
rect 6880 -1000 8880 -985
rect 9145 985 11145 1000
rect 9145 -985 9160 985
rect 11130 -985 11145 985
rect 9145 -1000 11145 -985
rect 11410 985 13410 1000
rect 11410 -985 11425 985
rect 13395 -985 13410 985
rect 11410 -1000 13410 -985
rect -13505 -1175 -11505 -1160
rect -13505 -3145 -13490 -1175
rect -11520 -3145 -11505 -1175
rect -13505 -3160 -11505 -3145
rect -11240 -1175 -9240 -1160
rect -11240 -3145 -11225 -1175
rect -9255 -3145 -9240 -1175
rect -11240 -3160 -9240 -3145
rect -8975 -1175 -6975 -1160
rect -8975 -3145 -8960 -1175
rect -6990 -3145 -6975 -1175
rect -8975 -3160 -6975 -3145
rect -6710 -1175 -4710 -1160
rect -6710 -3145 -6695 -1175
rect -4725 -3145 -4710 -1175
rect -6710 -3160 -4710 -3145
rect -4445 -1175 -2445 -1160
rect -4445 -3145 -4430 -1175
rect -2460 -3145 -2445 -1175
rect -4445 -3160 -2445 -3145
rect -2180 -1175 -180 -1160
rect -2180 -3145 -2165 -1175
rect -195 -3145 -180 -1175
rect -2180 -3160 -180 -3145
rect 85 -1175 2085 -1160
rect 85 -3145 100 -1175
rect 2070 -3145 2085 -1175
rect 85 -3160 2085 -3145
rect 2350 -1175 4350 -1160
rect 2350 -3145 2365 -1175
rect 4335 -3145 4350 -1175
rect 2350 -3160 4350 -3145
rect 4615 -1175 6615 -1160
rect 4615 -3145 4630 -1175
rect 6600 -3145 6615 -1175
rect 4615 -3160 6615 -3145
rect 6880 -1175 8880 -1160
rect 6880 -3145 6895 -1175
rect 8865 -3145 8880 -1175
rect 6880 -3160 8880 -3145
rect 9145 -1175 11145 -1160
rect 9145 -3145 9160 -1175
rect 11130 -3145 11145 -1175
rect 9145 -3160 11145 -3145
rect 11410 -1175 13410 -1160
rect 11410 -3145 11425 -1175
rect 13395 -3145 13410 -1175
rect 11410 -3160 13410 -3145
rect -13505 -3335 -11505 -3320
rect -13505 -5305 -13490 -3335
rect -11520 -5305 -11505 -3335
rect -13505 -5320 -11505 -5305
rect -11240 -3335 -9240 -3320
rect -11240 -5305 -11225 -3335
rect -9255 -5305 -9240 -3335
rect -11240 -5320 -9240 -5305
rect -8975 -3335 -6975 -3320
rect -8975 -5305 -8960 -3335
rect -6990 -5305 -6975 -3335
rect -8975 -5320 -6975 -5305
rect -6710 -3335 -4710 -3320
rect -6710 -5305 -6695 -3335
rect -4725 -5305 -4710 -3335
rect -6710 -5320 -4710 -5305
rect -4445 -3335 -2445 -3320
rect -4445 -5305 -4430 -3335
rect -2460 -5305 -2445 -3335
rect -4445 -5320 -2445 -5305
rect -2180 -3335 -180 -3320
rect -2180 -5305 -2165 -3335
rect -195 -5305 -180 -3335
rect -2180 -5320 -180 -5305
rect 85 -3335 2085 -3320
rect 85 -5305 100 -3335
rect 2070 -5305 2085 -3335
rect 85 -5320 2085 -5305
rect 2350 -3335 4350 -3320
rect 2350 -5305 2365 -3335
rect 4335 -5305 4350 -3335
rect 2350 -5320 4350 -5305
rect 4615 -3335 6615 -3320
rect 4615 -5305 4630 -3335
rect 6600 -5305 6615 -3335
rect 4615 -5320 6615 -5305
rect 6880 -3335 8880 -3320
rect 6880 -5305 6895 -3335
rect 8865 -5305 8880 -3335
rect 6880 -5320 8880 -5305
rect 9145 -3335 11145 -3320
rect 9145 -5305 9160 -3335
rect 11130 -5305 11145 -3335
rect 9145 -5320 11145 -5305
rect 11410 -3335 13410 -3320
rect 11410 -5305 11425 -3335
rect 13395 -5305 13410 -3335
rect 11410 -5320 13410 -5305
rect -13505 -5495 -11505 -5480
rect -13505 -7465 -13490 -5495
rect -11520 -7465 -11505 -5495
rect -13505 -7480 -11505 -7465
rect -11240 -5495 -9240 -5480
rect -11240 -7465 -11225 -5495
rect -9255 -7465 -9240 -5495
rect -11240 -7480 -9240 -7465
rect -8975 -5495 -6975 -5480
rect -8975 -7465 -8960 -5495
rect -6990 -7465 -6975 -5495
rect -8975 -7480 -6975 -7465
rect -6710 -5495 -4710 -5480
rect -6710 -7465 -6695 -5495
rect -4725 -7465 -4710 -5495
rect -6710 -7480 -4710 -7465
rect -4445 -5495 -2445 -5480
rect -4445 -7465 -4430 -5495
rect -2460 -7465 -2445 -5495
rect -4445 -7480 -2445 -7465
rect -2180 -5495 -180 -5480
rect -2180 -7465 -2165 -5495
rect -195 -7465 -180 -5495
rect -2180 -7480 -180 -7465
rect 85 -5495 2085 -5480
rect 85 -7465 100 -5495
rect 2070 -7465 2085 -5495
rect 85 -7480 2085 -7465
rect 2350 -5495 4350 -5480
rect 2350 -7465 2365 -5495
rect 4335 -7465 4350 -5495
rect 2350 -7480 4350 -7465
rect 4615 -5495 6615 -5480
rect 4615 -7465 4630 -5495
rect 6600 -7465 6615 -5495
rect 4615 -7480 6615 -7465
rect 6880 -5495 8880 -5480
rect 6880 -7465 6895 -5495
rect 8865 -7465 8880 -5495
rect 6880 -7480 8880 -7465
rect 9145 -5495 11145 -5480
rect 9145 -7465 9160 -5495
rect 11130 -7465 11145 -5495
rect 9145 -7480 11145 -7465
rect 11410 -5495 13410 -5480
rect 11410 -7465 11425 -5495
rect 13395 -7465 13410 -5495
rect 11410 -7480 13410 -7465
<< mimcapcontact >>
rect -13490 5495 -11520 7465
rect -11225 5495 -9255 7465
rect -8960 5495 -6990 7465
rect -6695 5495 -4725 7465
rect -4430 5495 -2460 7465
rect -2165 5495 -195 7465
rect 100 5495 2070 7465
rect 2365 5495 4335 7465
rect 4630 5495 6600 7465
rect 6895 5495 8865 7465
rect 9160 5495 11130 7465
rect 11425 5495 13395 7465
rect -13490 3335 -11520 5305
rect -11225 3335 -9255 5305
rect -8960 3335 -6990 5305
rect -6695 3335 -4725 5305
rect -4430 3335 -2460 5305
rect -2165 3335 -195 5305
rect 100 3335 2070 5305
rect 2365 3335 4335 5305
rect 4630 3335 6600 5305
rect 6895 3335 8865 5305
rect 9160 3335 11130 5305
rect 11425 3335 13395 5305
rect -13490 1175 -11520 3145
rect -11225 1175 -9255 3145
rect -8960 1175 -6990 3145
rect -6695 1175 -4725 3145
rect -4430 1175 -2460 3145
rect -2165 1175 -195 3145
rect 100 1175 2070 3145
rect 2365 1175 4335 3145
rect 4630 1175 6600 3145
rect 6895 1175 8865 3145
rect 9160 1175 11130 3145
rect 11425 1175 13395 3145
rect -13490 -985 -11520 985
rect -11225 -985 -9255 985
rect -8960 -985 -6990 985
rect -6695 -985 -4725 985
rect -4430 -985 -2460 985
rect -2165 -985 -195 985
rect 100 -985 2070 985
rect 2365 -985 4335 985
rect 4630 -985 6600 985
rect 6895 -985 8865 985
rect 9160 -985 11130 985
rect 11425 -985 13395 985
rect -13490 -3145 -11520 -1175
rect -11225 -3145 -9255 -1175
rect -8960 -3145 -6990 -1175
rect -6695 -3145 -4725 -1175
rect -4430 -3145 -2460 -1175
rect -2165 -3145 -195 -1175
rect 100 -3145 2070 -1175
rect 2365 -3145 4335 -1175
rect 4630 -3145 6600 -1175
rect 6895 -3145 8865 -1175
rect 9160 -3145 11130 -1175
rect 11425 -3145 13395 -1175
rect -13490 -5305 -11520 -3335
rect -11225 -5305 -9255 -3335
rect -8960 -5305 -6990 -3335
rect -6695 -5305 -4725 -3335
rect -4430 -5305 -2460 -3335
rect -2165 -5305 -195 -3335
rect 100 -5305 2070 -3335
rect 2365 -5305 4335 -3335
rect 4630 -5305 6600 -3335
rect 6895 -5305 8865 -3335
rect 9160 -5305 11130 -3335
rect 11425 -5305 13395 -3335
rect -13490 -7465 -11520 -5495
rect -11225 -7465 -9255 -5495
rect -8960 -7465 -6990 -5495
rect -6695 -7465 -4725 -5495
rect -4430 -7465 -2460 -5495
rect -2165 -7465 -195 -5495
rect 100 -7465 2070 -5495
rect 2365 -7465 4335 -5495
rect 4630 -7465 6600 -5495
rect 6895 -7465 8865 -5495
rect 9160 -7465 11130 -5495
rect 11425 -7465 13395 -5495
<< metal4 >>
rect -13555 7516 -11360 7530
rect -13555 7480 -11420 7516
rect -13555 5480 -13505 7480
rect -11505 5480 -11420 7480
rect -13555 5444 -11420 5480
rect -11370 5444 -11360 7516
rect -13555 5430 -11360 5444
rect -11290 7516 -9095 7530
rect -11290 7480 -9155 7516
rect -11290 5480 -11240 7480
rect -9240 5480 -9155 7480
rect -11290 5444 -9155 5480
rect -9105 5444 -9095 7516
rect -11290 5430 -9095 5444
rect -9025 7516 -6830 7530
rect -9025 7480 -6890 7516
rect -9025 5480 -8975 7480
rect -6975 5480 -6890 7480
rect -9025 5444 -6890 5480
rect -6840 5444 -6830 7516
rect -9025 5430 -6830 5444
rect -6760 7516 -4565 7530
rect -6760 7480 -4625 7516
rect -6760 5480 -6710 7480
rect -4710 5480 -4625 7480
rect -6760 5444 -4625 5480
rect -4575 5444 -4565 7516
rect -6760 5430 -4565 5444
rect -4495 7516 -2300 7530
rect -4495 7480 -2360 7516
rect -4495 5480 -4445 7480
rect -2445 5480 -2360 7480
rect -4495 5444 -2360 5480
rect -2310 5444 -2300 7516
rect -4495 5430 -2300 5444
rect -2230 7516 -35 7530
rect -2230 7480 -95 7516
rect -2230 5480 -2180 7480
rect -180 5480 -95 7480
rect -2230 5444 -95 5480
rect -45 5444 -35 7516
rect -2230 5430 -35 5444
rect 35 7516 2230 7530
rect 35 7480 2170 7516
rect 35 5480 85 7480
rect 2085 5480 2170 7480
rect 35 5444 2170 5480
rect 2220 5444 2230 7516
rect 35 5430 2230 5444
rect 2300 7516 4495 7530
rect 2300 7480 4435 7516
rect 2300 5480 2350 7480
rect 4350 5480 4435 7480
rect 2300 5444 4435 5480
rect 4485 5444 4495 7516
rect 2300 5430 4495 5444
rect 4565 7516 6760 7530
rect 4565 7480 6700 7516
rect 4565 5480 4615 7480
rect 6615 5480 6700 7480
rect 4565 5444 6700 5480
rect 6750 5444 6760 7516
rect 4565 5430 6760 5444
rect 6830 7516 9025 7530
rect 6830 7480 8965 7516
rect 6830 5480 6880 7480
rect 8880 5480 8965 7480
rect 6830 5444 8965 5480
rect 9015 5444 9025 7516
rect 6830 5430 9025 5444
rect 9095 7516 11290 7530
rect 9095 7480 11230 7516
rect 9095 5480 9145 7480
rect 11145 5480 11230 7480
rect 9095 5444 11230 5480
rect 11280 5444 11290 7516
rect 9095 5430 11290 5444
rect 11360 7516 13555 7530
rect 11360 7480 13495 7516
rect 11360 5480 11410 7480
rect 13410 5480 13495 7480
rect 11360 5444 13495 5480
rect 13545 5444 13555 7516
rect 11360 5430 13555 5444
rect -13555 5356 -11360 5370
rect -13555 5320 -11420 5356
rect -13555 3320 -13505 5320
rect -11505 3320 -11420 5320
rect -13555 3284 -11420 3320
rect -11370 3284 -11360 5356
rect -13555 3270 -11360 3284
rect -11290 5356 -9095 5370
rect -11290 5320 -9155 5356
rect -11290 3320 -11240 5320
rect -9240 3320 -9155 5320
rect -11290 3284 -9155 3320
rect -9105 3284 -9095 5356
rect -11290 3270 -9095 3284
rect -9025 5356 -6830 5370
rect -9025 5320 -6890 5356
rect -9025 3320 -8975 5320
rect -6975 3320 -6890 5320
rect -9025 3284 -6890 3320
rect -6840 3284 -6830 5356
rect -9025 3270 -6830 3284
rect -6760 5356 -4565 5370
rect -6760 5320 -4625 5356
rect -6760 3320 -6710 5320
rect -4710 3320 -4625 5320
rect -6760 3284 -4625 3320
rect -4575 3284 -4565 5356
rect -6760 3270 -4565 3284
rect -4495 5356 -2300 5370
rect -4495 5320 -2360 5356
rect -4495 3320 -4445 5320
rect -2445 3320 -2360 5320
rect -4495 3284 -2360 3320
rect -2310 3284 -2300 5356
rect -4495 3270 -2300 3284
rect -2230 5356 -35 5370
rect -2230 5320 -95 5356
rect -2230 3320 -2180 5320
rect -180 3320 -95 5320
rect -2230 3284 -95 3320
rect -45 3284 -35 5356
rect -2230 3270 -35 3284
rect 35 5356 2230 5370
rect 35 5320 2170 5356
rect 35 3320 85 5320
rect 2085 3320 2170 5320
rect 35 3284 2170 3320
rect 2220 3284 2230 5356
rect 35 3270 2230 3284
rect 2300 5356 4495 5370
rect 2300 5320 4435 5356
rect 2300 3320 2350 5320
rect 4350 3320 4435 5320
rect 2300 3284 4435 3320
rect 4485 3284 4495 5356
rect 2300 3270 4495 3284
rect 4565 5356 6760 5370
rect 4565 5320 6700 5356
rect 4565 3320 4615 5320
rect 6615 3320 6700 5320
rect 4565 3284 6700 3320
rect 6750 3284 6760 5356
rect 4565 3270 6760 3284
rect 6830 5356 9025 5370
rect 6830 5320 8965 5356
rect 6830 3320 6880 5320
rect 8880 3320 8965 5320
rect 6830 3284 8965 3320
rect 9015 3284 9025 5356
rect 6830 3270 9025 3284
rect 9095 5356 11290 5370
rect 9095 5320 11230 5356
rect 9095 3320 9145 5320
rect 11145 3320 11230 5320
rect 9095 3284 11230 3320
rect 11280 3284 11290 5356
rect 9095 3270 11290 3284
rect 11360 5356 13555 5370
rect 11360 5320 13495 5356
rect 11360 3320 11410 5320
rect 13410 3320 13495 5320
rect 11360 3284 13495 3320
rect 13545 3284 13555 5356
rect 11360 3270 13555 3284
rect -13555 3196 -11360 3210
rect -13555 3160 -11420 3196
rect -13555 1160 -13505 3160
rect -11505 1160 -11420 3160
rect -13555 1124 -11420 1160
rect -11370 1124 -11360 3196
rect -13555 1110 -11360 1124
rect -11290 3196 -9095 3210
rect -11290 3160 -9155 3196
rect -11290 1160 -11240 3160
rect -9240 1160 -9155 3160
rect -11290 1124 -9155 1160
rect -9105 1124 -9095 3196
rect -11290 1110 -9095 1124
rect -9025 3196 -6830 3210
rect -9025 3160 -6890 3196
rect -9025 1160 -8975 3160
rect -6975 1160 -6890 3160
rect -9025 1124 -6890 1160
rect -6840 1124 -6830 3196
rect -9025 1110 -6830 1124
rect -6760 3196 -4565 3210
rect -6760 3160 -4625 3196
rect -6760 1160 -6710 3160
rect -4710 1160 -4625 3160
rect -6760 1124 -4625 1160
rect -4575 1124 -4565 3196
rect -6760 1110 -4565 1124
rect -4495 3196 -2300 3210
rect -4495 3160 -2360 3196
rect -4495 1160 -4445 3160
rect -2445 1160 -2360 3160
rect -4495 1124 -2360 1160
rect -2310 1124 -2300 3196
rect -4495 1110 -2300 1124
rect -2230 3196 -35 3210
rect -2230 3160 -95 3196
rect -2230 1160 -2180 3160
rect -180 1160 -95 3160
rect -2230 1124 -95 1160
rect -45 1124 -35 3196
rect -2230 1110 -35 1124
rect 35 3196 2230 3210
rect 35 3160 2170 3196
rect 35 1160 85 3160
rect 2085 1160 2170 3160
rect 35 1124 2170 1160
rect 2220 1124 2230 3196
rect 35 1110 2230 1124
rect 2300 3196 4495 3210
rect 2300 3160 4435 3196
rect 2300 1160 2350 3160
rect 4350 1160 4435 3160
rect 2300 1124 4435 1160
rect 4485 1124 4495 3196
rect 2300 1110 4495 1124
rect 4565 3196 6760 3210
rect 4565 3160 6700 3196
rect 4565 1160 4615 3160
rect 6615 1160 6700 3160
rect 4565 1124 6700 1160
rect 6750 1124 6760 3196
rect 4565 1110 6760 1124
rect 6830 3196 9025 3210
rect 6830 3160 8965 3196
rect 6830 1160 6880 3160
rect 8880 1160 8965 3160
rect 6830 1124 8965 1160
rect 9015 1124 9025 3196
rect 6830 1110 9025 1124
rect 9095 3196 11290 3210
rect 9095 3160 11230 3196
rect 9095 1160 9145 3160
rect 11145 1160 11230 3160
rect 9095 1124 11230 1160
rect 11280 1124 11290 3196
rect 9095 1110 11290 1124
rect 11360 3196 13555 3210
rect 11360 3160 13495 3196
rect 11360 1160 11410 3160
rect 13410 1160 13495 3160
rect 11360 1124 13495 1160
rect 13545 1124 13555 3196
rect 11360 1110 13555 1124
rect -13555 1036 -11360 1050
rect -13555 1000 -11420 1036
rect -13555 -1000 -13505 1000
rect -11505 -1000 -11420 1000
rect -13555 -1036 -11420 -1000
rect -11370 -1036 -11360 1036
rect -13555 -1050 -11360 -1036
rect -11290 1036 -9095 1050
rect -11290 1000 -9155 1036
rect -11290 -1000 -11240 1000
rect -9240 -1000 -9155 1000
rect -11290 -1036 -9155 -1000
rect -9105 -1036 -9095 1036
rect -11290 -1050 -9095 -1036
rect -9025 1036 -6830 1050
rect -9025 1000 -6890 1036
rect -9025 -1000 -8975 1000
rect -6975 -1000 -6890 1000
rect -9025 -1036 -6890 -1000
rect -6840 -1036 -6830 1036
rect -9025 -1050 -6830 -1036
rect -6760 1036 -4565 1050
rect -6760 1000 -4625 1036
rect -6760 -1000 -6710 1000
rect -4710 -1000 -4625 1000
rect -6760 -1036 -4625 -1000
rect -4575 -1036 -4565 1036
rect -6760 -1050 -4565 -1036
rect -4495 1036 -2300 1050
rect -4495 1000 -2360 1036
rect -4495 -1000 -4445 1000
rect -2445 -1000 -2360 1000
rect -4495 -1036 -2360 -1000
rect -2310 -1036 -2300 1036
rect -4495 -1050 -2300 -1036
rect -2230 1036 -35 1050
rect -2230 1000 -95 1036
rect -2230 -1000 -2180 1000
rect -180 -1000 -95 1000
rect -2230 -1036 -95 -1000
rect -45 -1036 -35 1036
rect -2230 -1050 -35 -1036
rect 35 1036 2230 1050
rect 35 1000 2170 1036
rect 35 -1000 85 1000
rect 2085 -1000 2170 1000
rect 35 -1036 2170 -1000
rect 2220 -1036 2230 1036
rect 35 -1050 2230 -1036
rect 2300 1036 4495 1050
rect 2300 1000 4435 1036
rect 2300 -1000 2350 1000
rect 4350 -1000 4435 1000
rect 2300 -1036 4435 -1000
rect 4485 -1036 4495 1036
rect 2300 -1050 4495 -1036
rect 4565 1036 6760 1050
rect 4565 1000 6700 1036
rect 4565 -1000 4615 1000
rect 6615 -1000 6700 1000
rect 4565 -1036 6700 -1000
rect 6750 -1036 6760 1036
rect 4565 -1050 6760 -1036
rect 6830 1036 9025 1050
rect 6830 1000 8965 1036
rect 6830 -1000 6880 1000
rect 8880 -1000 8965 1000
rect 6830 -1036 8965 -1000
rect 9015 -1036 9025 1036
rect 6830 -1050 9025 -1036
rect 9095 1036 11290 1050
rect 9095 1000 11230 1036
rect 9095 -1000 9145 1000
rect 11145 -1000 11230 1000
rect 9095 -1036 11230 -1000
rect 11280 -1036 11290 1036
rect 9095 -1050 11290 -1036
rect 11360 1036 13555 1050
rect 11360 1000 13495 1036
rect 11360 -1000 11410 1000
rect 13410 -1000 13495 1000
rect 11360 -1036 13495 -1000
rect 13545 -1036 13555 1036
rect 11360 -1050 13555 -1036
rect -13555 -1124 -11360 -1110
rect -13555 -1160 -11420 -1124
rect -13555 -3160 -13505 -1160
rect -11505 -3160 -11420 -1160
rect -13555 -3196 -11420 -3160
rect -11370 -3196 -11360 -1124
rect -13555 -3210 -11360 -3196
rect -11290 -1124 -9095 -1110
rect -11290 -1160 -9155 -1124
rect -11290 -3160 -11240 -1160
rect -9240 -3160 -9155 -1160
rect -11290 -3196 -9155 -3160
rect -9105 -3196 -9095 -1124
rect -11290 -3210 -9095 -3196
rect -9025 -1124 -6830 -1110
rect -9025 -1160 -6890 -1124
rect -9025 -3160 -8975 -1160
rect -6975 -3160 -6890 -1160
rect -9025 -3196 -6890 -3160
rect -6840 -3196 -6830 -1124
rect -9025 -3210 -6830 -3196
rect -6760 -1124 -4565 -1110
rect -6760 -1160 -4625 -1124
rect -6760 -3160 -6710 -1160
rect -4710 -3160 -4625 -1160
rect -6760 -3196 -4625 -3160
rect -4575 -3196 -4565 -1124
rect -6760 -3210 -4565 -3196
rect -4495 -1124 -2300 -1110
rect -4495 -1160 -2360 -1124
rect -4495 -3160 -4445 -1160
rect -2445 -3160 -2360 -1160
rect -4495 -3196 -2360 -3160
rect -2310 -3196 -2300 -1124
rect -4495 -3210 -2300 -3196
rect -2230 -1124 -35 -1110
rect -2230 -1160 -95 -1124
rect -2230 -3160 -2180 -1160
rect -180 -3160 -95 -1160
rect -2230 -3196 -95 -3160
rect -45 -3196 -35 -1124
rect -2230 -3210 -35 -3196
rect 35 -1124 2230 -1110
rect 35 -1160 2170 -1124
rect 35 -3160 85 -1160
rect 2085 -3160 2170 -1160
rect 35 -3196 2170 -3160
rect 2220 -3196 2230 -1124
rect 35 -3210 2230 -3196
rect 2300 -1124 4495 -1110
rect 2300 -1160 4435 -1124
rect 2300 -3160 2350 -1160
rect 4350 -3160 4435 -1160
rect 2300 -3196 4435 -3160
rect 4485 -3196 4495 -1124
rect 2300 -3210 4495 -3196
rect 4565 -1124 6760 -1110
rect 4565 -1160 6700 -1124
rect 4565 -3160 4615 -1160
rect 6615 -3160 6700 -1160
rect 4565 -3196 6700 -3160
rect 6750 -3196 6760 -1124
rect 4565 -3210 6760 -3196
rect 6830 -1124 9025 -1110
rect 6830 -1160 8965 -1124
rect 6830 -3160 6880 -1160
rect 8880 -3160 8965 -1160
rect 6830 -3196 8965 -3160
rect 9015 -3196 9025 -1124
rect 6830 -3210 9025 -3196
rect 9095 -1124 11290 -1110
rect 9095 -1160 11230 -1124
rect 9095 -3160 9145 -1160
rect 11145 -3160 11230 -1160
rect 9095 -3196 11230 -3160
rect 11280 -3196 11290 -1124
rect 9095 -3210 11290 -3196
rect 11360 -1124 13555 -1110
rect 11360 -1160 13495 -1124
rect 11360 -3160 11410 -1160
rect 13410 -3160 13495 -1160
rect 11360 -3196 13495 -3160
rect 13545 -3196 13555 -1124
rect 11360 -3210 13555 -3196
rect -13555 -3284 -11360 -3270
rect -13555 -3320 -11420 -3284
rect -13555 -5320 -13505 -3320
rect -11505 -5320 -11420 -3320
rect -13555 -5356 -11420 -5320
rect -11370 -5356 -11360 -3284
rect -13555 -5370 -11360 -5356
rect -11290 -3284 -9095 -3270
rect -11290 -3320 -9155 -3284
rect -11290 -5320 -11240 -3320
rect -9240 -5320 -9155 -3320
rect -11290 -5356 -9155 -5320
rect -9105 -5356 -9095 -3284
rect -11290 -5370 -9095 -5356
rect -9025 -3284 -6830 -3270
rect -9025 -3320 -6890 -3284
rect -9025 -5320 -8975 -3320
rect -6975 -5320 -6890 -3320
rect -9025 -5356 -6890 -5320
rect -6840 -5356 -6830 -3284
rect -9025 -5370 -6830 -5356
rect -6760 -3284 -4565 -3270
rect -6760 -3320 -4625 -3284
rect -6760 -5320 -6710 -3320
rect -4710 -5320 -4625 -3320
rect -6760 -5356 -4625 -5320
rect -4575 -5356 -4565 -3284
rect -6760 -5370 -4565 -5356
rect -4495 -3284 -2300 -3270
rect -4495 -3320 -2360 -3284
rect -4495 -5320 -4445 -3320
rect -2445 -5320 -2360 -3320
rect -4495 -5356 -2360 -5320
rect -2310 -5356 -2300 -3284
rect -4495 -5370 -2300 -5356
rect -2230 -3284 -35 -3270
rect -2230 -3320 -95 -3284
rect -2230 -5320 -2180 -3320
rect -180 -5320 -95 -3320
rect -2230 -5356 -95 -5320
rect -45 -5356 -35 -3284
rect -2230 -5370 -35 -5356
rect 35 -3284 2230 -3270
rect 35 -3320 2170 -3284
rect 35 -5320 85 -3320
rect 2085 -5320 2170 -3320
rect 35 -5356 2170 -5320
rect 2220 -5356 2230 -3284
rect 35 -5370 2230 -5356
rect 2300 -3284 4495 -3270
rect 2300 -3320 4435 -3284
rect 2300 -5320 2350 -3320
rect 4350 -5320 4435 -3320
rect 2300 -5356 4435 -5320
rect 4485 -5356 4495 -3284
rect 2300 -5370 4495 -5356
rect 4565 -3284 6760 -3270
rect 4565 -3320 6700 -3284
rect 4565 -5320 4615 -3320
rect 6615 -5320 6700 -3320
rect 4565 -5356 6700 -5320
rect 6750 -5356 6760 -3284
rect 4565 -5370 6760 -5356
rect 6830 -3284 9025 -3270
rect 6830 -3320 8965 -3284
rect 6830 -5320 6880 -3320
rect 8880 -5320 8965 -3320
rect 6830 -5356 8965 -5320
rect 9015 -5356 9025 -3284
rect 6830 -5370 9025 -5356
rect 9095 -3284 11290 -3270
rect 9095 -3320 11230 -3284
rect 9095 -5320 9145 -3320
rect 11145 -5320 11230 -3320
rect 9095 -5356 11230 -5320
rect 11280 -5356 11290 -3284
rect 9095 -5370 11290 -5356
rect 11360 -3284 13555 -3270
rect 11360 -3320 13495 -3284
rect 11360 -5320 11410 -3320
rect 13410 -5320 13495 -3320
rect 11360 -5356 13495 -5320
rect 13545 -5356 13555 -3284
rect 11360 -5370 13555 -5356
rect -13555 -5444 -11360 -5430
rect -13555 -5480 -11420 -5444
rect -13555 -7480 -13505 -5480
rect -11505 -7480 -11420 -5480
rect -13555 -7516 -11420 -7480
rect -11370 -7516 -11360 -5444
rect -13555 -7530 -11360 -7516
rect -11290 -5444 -9095 -5430
rect -11290 -5480 -9155 -5444
rect -11290 -7480 -11240 -5480
rect -9240 -7480 -9155 -5480
rect -11290 -7516 -9155 -7480
rect -9105 -7516 -9095 -5444
rect -11290 -7530 -9095 -7516
rect -9025 -5444 -6830 -5430
rect -9025 -5480 -6890 -5444
rect -9025 -7480 -8975 -5480
rect -6975 -7480 -6890 -5480
rect -9025 -7516 -6890 -7480
rect -6840 -7516 -6830 -5444
rect -9025 -7530 -6830 -7516
rect -6760 -5444 -4565 -5430
rect -6760 -5480 -4625 -5444
rect -6760 -7480 -6710 -5480
rect -4710 -7480 -4625 -5480
rect -6760 -7516 -4625 -7480
rect -4575 -7516 -4565 -5444
rect -6760 -7530 -4565 -7516
rect -4495 -5444 -2300 -5430
rect -4495 -5480 -2360 -5444
rect -4495 -7480 -4445 -5480
rect -2445 -7480 -2360 -5480
rect -4495 -7516 -2360 -7480
rect -2310 -7516 -2300 -5444
rect -4495 -7530 -2300 -7516
rect -2230 -5444 -35 -5430
rect -2230 -5480 -95 -5444
rect -2230 -7480 -2180 -5480
rect -180 -7480 -95 -5480
rect -2230 -7516 -95 -7480
rect -45 -7516 -35 -5444
rect -2230 -7530 -35 -7516
rect 35 -5444 2230 -5430
rect 35 -5480 2170 -5444
rect 35 -7480 85 -5480
rect 2085 -7480 2170 -5480
rect 35 -7516 2170 -7480
rect 2220 -7516 2230 -5444
rect 35 -7530 2230 -7516
rect 2300 -5444 4495 -5430
rect 2300 -5480 4435 -5444
rect 2300 -7480 2350 -5480
rect 4350 -7480 4435 -5480
rect 2300 -7516 4435 -7480
rect 4485 -7516 4495 -5444
rect 2300 -7530 4495 -7516
rect 4565 -5444 6760 -5430
rect 4565 -5480 6700 -5444
rect 4565 -7480 4615 -5480
rect 6615 -7480 6700 -5480
rect 4565 -7516 6700 -7480
rect 6750 -7516 6760 -5444
rect 4565 -7530 6760 -7516
rect 6830 -5444 9025 -5430
rect 6830 -5480 8965 -5444
rect 6830 -7480 6880 -5480
rect 8880 -7480 8965 -5480
rect 6830 -7516 8965 -7480
rect 9015 -7516 9025 -5444
rect 6830 -7530 9025 -7516
rect 9095 -5444 11290 -5430
rect 9095 -5480 11230 -5444
rect 9095 -7480 9145 -5480
rect 11145 -7480 11230 -5480
rect 9095 -7516 11230 -7480
rect 11280 -7516 11290 -5444
rect 9095 -7530 11290 -7516
rect 11360 -5444 13555 -5430
rect 11360 -5480 13495 -5444
rect 11360 -7480 11410 -5480
rect 13410 -7480 13495 -5480
rect 11360 -7516 13495 -7480
rect 13545 -7516 13555 -5444
rect 11360 -7530 13555 -7516
<< viatp >>
rect -11420 5444 -11370 7516
rect -9155 5444 -9105 7516
rect -6890 5444 -6840 7516
rect -4625 5444 -4575 7516
rect -2360 5444 -2310 7516
rect -95 5444 -45 7516
rect 2170 5444 2220 7516
rect 4435 5444 4485 7516
rect 6700 5444 6750 7516
rect 8965 5444 9015 7516
rect 11230 5444 11280 7516
rect 13495 5444 13545 7516
rect -11420 3284 -11370 5356
rect -9155 3284 -9105 5356
rect -6890 3284 -6840 5356
rect -4625 3284 -4575 5356
rect -2360 3284 -2310 5356
rect -95 3284 -45 5356
rect 2170 3284 2220 5356
rect 4435 3284 4485 5356
rect 6700 3284 6750 5356
rect 8965 3284 9015 5356
rect 11230 3284 11280 5356
rect 13495 3284 13545 5356
rect -11420 1124 -11370 3196
rect -9155 1124 -9105 3196
rect -6890 1124 -6840 3196
rect -4625 1124 -4575 3196
rect -2360 1124 -2310 3196
rect -95 1124 -45 3196
rect 2170 1124 2220 3196
rect 4435 1124 4485 3196
rect 6700 1124 6750 3196
rect 8965 1124 9015 3196
rect 11230 1124 11280 3196
rect 13495 1124 13545 3196
rect -11420 -1036 -11370 1036
rect -9155 -1036 -9105 1036
rect -6890 -1036 -6840 1036
rect -4625 -1036 -4575 1036
rect -2360 -1036 -2310 1036
rect -95 -1036 -45 1036
rect 2170 -1036 2220 1036
rect 4435 -1036 4485 1036
rect 6700 -1036 6750 1036
rect 8965 -1036 9015 1036
rect 11230 -1036 11280 1036
rect 13495 -1036 13545 1036
rect -11420 -3196 -11370 -1124
rect -9155 -3196 -9105 -1124
rect -6890 -3196 -6840 -1124
rect -4625 -3196 -4575 -1124
rect -2360 -3196 -2310 -1124
rect -95 -3196 -45 -1124
rect 2170 -3196 2220 -1124
rect 4435 -3196 4485 -1124
rect 6700 -3196 6750 -1124
rect 8965 -3196 9015 -1124
rect 11230 -3196 11280 -1124
rect 13495 -3196 13545 -1124
rect -11420 -5356 -11370 -3284
rect -9155 -5356 -9105 -3284
rect -6890 -5356 -6840 -3284
rect -4625 -5356 -4575 -3284
rect -2360 -5356 -2310 -3284
rect -95 -5356 -45 -3284
rect 2170 -5356 2220 -3284
rect 4435 -5356 4485 -3284
rect 6700 -5356 6750 -3284
rect 8965 -5356 9015 -3284
rect 11230 -5356 11280 -3284
rect 13495 -5356 13545 -3284
rect -11420 -7516 -11370 -5444
rect -9155 -7516 -9105 -5444
rect -6890 -7516 -6840 -5444
rect -4625 -7516 -4575 -5444
rect -2360 -7516 -2310 -5444
rect -95 -7516 -45 -5444
rect 2170 -7516 2220 -5444
rect 4435 -7516 4485 -5444
rect 6700 -7516 6750 -5444
rect 8965 -7516 9015 -5444
rect 11230 -7516 11280 -5444
rect 13495 -7516 13545 -5444
<< metaltp >>
rect -12540 7465 -12470 7560
rect -11430 7516 -11360 7560
rect -12540 5305 -12470 5495
rect -11430 5444 -11420 7516
rect -11370 5444 -11360 7516
rect -10275 7465 -10205 7560
rect -9165 7516 -9095 7560
rect -11430 5356 -11360 5444
rect -12540 3145 -12470 3335
rect -11430 3284 -11420 5356
rect -11370 3284 -11360 5356
rect -10275 5305 -10205 5495
rect -9165 5444 -9155 7516
rect -9105 5444 -9095 7516
rect -8010 7465 -7940 7560
rect -6900 7516 -6830 7560
rect -9165 5356 -9095 5444
rect -11430 3196 -11360 3284
rect -12540 985 -12470 1175
rect -11430 1124 -11420 3196
rect -11370 1124 -11360 3196
rect -10275 3145 -10205 3335
rect -9165 3284 -9155 5356
rect -9105 3284 -9095 5356
rect -8010 5305 -7940 5495
rect -6900 5444 -6890 7516
rect -6840 5444 -6830 7516
rect -5745 7465 -5675 7560
rect -4635 7516 -4565 7560
rect -6900 5356 -6830 5444
rect -9165 3196 -9095 3284
rect -11430 1036 -11360 1124
rect -12540 -1175 -12470 -985
rect -11430 -1036 -11420 1036
rect -11370 -1036 -11360 1036
rect -10275 985 -10205 1175
rect -9165 1124 -9155 3196
rect -9105 1124 -9095 3196
rect -8010 3145 -7940 3335
rect -6900 3284 -6890 5356
rect -6840 3284 -6830 5356
rect -5745 5305 -5675 5495
rect -4635 5444 -4625 7516
rect -4575 5444 -4565 7516
rect -3480 7465 -3410 7560
rect -2370 7516 -2300 7560
rect -4635 5356 -4565 5444
rect -6900 3196 -6830 3284
rect -9165 1036 -9095 1124
rect -11430 -1124 -11360 -1036
rect -12540 -3335 -12470 -3145
rect -11430 -3196 -11420 -1124
rect -11370 -3196 -11360 -1124
rect -10275 -1175 -10205 -985
rect -9165 -1036 -9155 1036
rect -9105 -1036 -9095 1036
rect -8010 985 -7940 1175
rect -6900 1124 -6890 3196
rect -6840 1124 -6830 3196
rect -5745 3145 -5675 3335
rect -4635 3284 -4625 5356
rect -4575 3284 -4565 5356
rect -3480 5305 -3410 5495
rect -2370 5444 -2360 7516
rect -2310 5444 -2300 7516
rect -1215 7465 -1145 7560
rect -105 7516 -35 7560
rect -2370 5356 -2300 5444
rect -4635 3196 -4565 3284
rect -6900 1036 -6830 1124
rect -9165 -1124 -9095 -1036
rect -11430 -3284 -11360 -3196
rect -12540 -5495 -12470 -5305
rect -11430 -5356 -11420 -3284
rect -11370 -5356 -11360 -3284
rect -10275 -3335 -10205 -3145
rect -9165 -3196 -9155 -1124
rect -9105 -3196 -9095 -1124
rect -8010 -1175 -7940 -985
rect -6900 -1036 -6890 1036
rect -6840 -1036 -6830 1036
rect -5745 985 -5675 1175
rect -4635 1124 -4625 3196
rect -4575 1124 -4565 3196
rect -3480 3145 -3410 3335
rect -2370 3284 -2360 5356
rect -2310 3284 -2300 5356
rect -1215 5305 -1145 5495
rect -105 5444 -95 7516
rect -45 5444 -35 7516
rect 1050 7465 1120 7560
rect 2160 7516 2230 7560
rect -105 5356 -35 5444
rect -2370 3196 -2300 3284
rect -4635 1036 -4565 1124
rect -6900 -1124 -6830 -1036
rect -9165 -3284 -9095 -3196
rect -11430 -5444 -11360 -5356
rect -12540 -7560 -12470 -7465
rect -11430 -7516 -11420 -5444
rect -11370 -7516 -11360 -5444
rect -10275 -5495 -10205 -5305
rect -9165 -5356 -9155 -3284
rect -9105 -5356 -9095 -3284
rect -8010 -3335 -7940 -3145
rect -6900 -3196 -6890 -1124
rect -6840 -3196 -6830 -1124
rect -5745 -1175 -5675 -985
rect -4635 -1036 -4625 1036
rect -4575 -1036 -4565 1036
rect -3480 985 -3410 1175
rect -2370 1124 -2360 3196
rect -2310 1124 -2300 3196
rect -1215 3145 -1145 3335
rect -105 3284 -95 5356
rect -45 3284 -35 5356
rect 1050 5305 1120 5495
rect 2160 5444 2170 7516
rect 2220 5444 2230 7516
rect 3315 7465 3385 7560
rect 4425 7516 4495 7560
rect 2160 5356 2230 5444
rect -105 3196 -35 3284
rect -2370 1036 -2300 1124
rect -4635 -1124 -4565 -1036
rect -6900 -3284 -6830 -3196
rect -9165 -5444 -9095 -5356
rect -11430 -7560 -11360 -7516
rect -10275 -7560 -10205 -7465
rect -9165 -7516 -9155 -5444
rect -9105 -7516 -9095 -5444
rect -8010 -5495 -7940 -5305
rect -6900 -5356 -6890 -3284
rect -6840 -5356 -6830 -3284
rect -5745 -3335 -5675 -3145
rect -4635 -3196 -4625 -1124
rect -4575 -3196 -4565 -1124
rect -3480 -1175 -3410 -985
rect -2370 -1036 -2360 1036
rect -2310 -1036 -2300 1036
rect -1215 985 -1145 1175
rect -105 1124 -95 3196
rect -45 1124 -35 3196
rect 1050 3145 1120 3335
rect 2160 3284 2170 5356
rect 2220 3284 2230 5356
rect 3315 5305 3385 5495
rect 4425 5444 4435 7516
rect 4485 5444 4495 7516
rect 5580 7465 5650 7560
rect 6690 7516 6760 7560
rect 4425 5356 4495 5444
rect 2160 3196 2230 3284
rect -105 1036 -35 1124
rect -2370 -1124 -2300 -1036
rect -4635 -3284 -4565 -3196
rect -6900 -5444 -6830 -5356
rect -9165 -7560 -9095 -7516
rect -8010 -7560 -7940 -7465
rect -6900 -7516 -6890 -5444
rect -6840 -7516 -6830 -5444
rect -5745 -5495 -5675 -5305
rect -4635 -5356 -4625 -3284
rect -4575 -5356 -4565 -3284
rect -3480 -3335 -3410 -3145
rect -2370 -3196 -2360 -1124
rect -2310 -3196 -2300 -1124
rect -1215 -1175 -1145 -985
rect -105 -1036 -95 1036
rect -45 -1036 -35 1036
rect 1050 985 1120 1175
rect 2160 1124 2170 3196
rect 2220 1124 2230 3196
rect 3315 3145 3385 3335
rect 4425 3284 4435 5356
rect 4485 3284 4495 5356
rect 5580 5305 5650 5495
rect 6690 5444 6700 7516
rect 6750 5444 6760 7516
rect 7845 7465 7915 7560
rect 8955 7516 9025 7560
rect 6690 5356 6760 5444
rect 4425 3196 4495 3284
rect 2160 1036 2230 1124
rect -105 -1124 -35 -1036
rect -2370 -3284 -2300 -3196
rect -4635 -5444 -4565 -5356
rect -6900 -7560 -6830 -7516
rect -5745 -7560 -5675 -7465
rect -4635 -7516 -4625 -5444
rect -4575 -7516 -4565 -5444
rect -3480 -5495 -3410 -5305
rect -2370 -5356 -2360 -3284
rect -2310 -5356 -2300 -3284
rect -1215 -3335 -1145 -3145
rect -105 -3196 -95 -1124
rect -45 -3196 -35 -1124
rect 1050 -1175 1120 -985
rect 2160 -1036 2170 1036
rect 2220 -1036 2230 1036
rect 3315 985 3385 1175
rect 4425 1124 4435 3196
rect 4485 1124 4495 3196
rect 5580 3145 5650 3335
rect 6690 3284 6700 5356
rect 6750 3284 6760 5356
rect 7845 5305 7915 5495
rect 8955 5444 8965 7516
rect 9015 5444 9025 7516
rect 10110 7465 10180 7560
rect 11220 7516 11290 7560
rect 8955 5356 9025 5444
rect 6690 3196 6760 3284
rect 4425 1036 4495 1124
rect 2160 -1124 2230 -1036
rect -105 -3284 -35 -3196
rect -2370 -5444 -2300 -5356
rect -4635 -7560 -4565 -7516
rect -3480 -7560 -3410 -7465
rect -2370 -7516 -2360 -5444
rect -2310 -7516 -2300 -5444
rect -1215 -5495 -1145 -5305
rect -105 -5356 -95 -3284
rect -45 -5356 -35 -3284
rect 1050 -3335 1120 -3145
rect 2160 -3196 2170 -1124
rect 2220 -3196 2230 -1124
rect 3315 -1175 3385 -985
rect 4425 -1036 4435 1036
rect 4485 -1036 4495 1036
rect 5580 985 5650 1175
rect 6690 1124 6700 3196
rect 6750 1124 6760 3196
rect 7845 3145 7915 3335
rect 8955 3284 8965 5356
rect 9015 3284 9025 5356
rect 10110 5305 10180 5495
rect 11220 5444 11230 7516
rect 11280 5444 11290 7516
rect 12375 7465 12445 7560
rect 13485 7516 13555 7560
rect 11220 5356 11290 5444
rect 8955 3196 9025 3284
rect 6690 1036 6760 1124
rect 4425 -1124 4495 -1036
rect 2160 -3284 2230 -3196
rect -105 -5444 -35 -5356
rect -2370 -7560 -2300 -7516
rect -1215 -7560 -1145 -7465
rect -105 -7516 -95 -5444
rect -45 -7516 -35 -5444
rect 1050 -5495 1120 -5305
rect 2160 -5356 2170 -3284
rect 2220 -5356 2230 -3284
rect 3315 -3335 3385 -3145
rect 4425 -3196 4435 -1124
rect 4485 -3196 4495 -1124
rect 5580 -1175 5650 -985
rect 6690 -1036 6700 1036
rect 6750 -1036 6760 1036
rect 7845 985 7915 1175
rect 8955 1124 8965 3196
rect 9015 1124 9025 3196
rect 10110 3145 10180 3335
rect 11220 3284 11230 5356
rect 11280 3284 11290 5356
rect 12375 5305 12445 5495
rect 13485 5444 13495 7516
rect 13545 5444 13555 7516
rect 13485 5356 13555 5444
rect 11220 3196 11290 3284
rect 8955 1036 9025 1124
rect 6690 -1124 6760 -1036
rect 4425 -3284 4495 -3196
rect 2160 -5444 2230 -5356
rect -105 -7560 -35 -7516
rect 1050 -7560 1120 -7465
rect 2160 -7516 2170 -5444
rect 2220 -7516 2230 -5444
rect 3315 -5495 3385 -5305
rect 4425 -5356 4435 -3284
rect 4485 -5356 4495 -3284
rect 5580 -3335 5650 -3145
rect 6690 -3196 6700 -1124
rect 6750 -3196 6760 -1124
rect 7845 -1175 7915 -985
rect 8955 -1036 8965 1036
rect 9015 -1036 9025 1036
rect 10110 985 10180 1175
rect 11220 1124 11230 3196
rect 11280 1124 11290 3196
rect 12375 3145 12445 3335
rect 13485 3284 13495 5356
rect 13545 3284 13555 5356
rect 13485 3196 13555 3284
rect 11220 1036 11290 1124
rect 8955 -1124 9025 -1036
rect 6690 -3284 6760 -3196
rect 4425 -5444 4495 -5356
rect 2160 -7560 2230 -7516
rect 3315 -7560 3385 -7465
rect 4425 -7516 4435 -5444
rect 4485 -7516 4495 -5444
rect 5580 -5495 5650 -5305
rect 6690 -5356 6700 -3284
rect 6750 -5356 6760 -3284
rect 7845 -3335 7915 -3145
rect 8955 -3196 8965 -1124
rect 9015 -3196 9025 -1124
rect 10110 -1175 10180 -985
rect 11220 -1036 11230 1036
rect 11280 -1036 11290 1036
rect 12375 985 12445 1175
rect 13485 1124 13495 3196
rect 13545 1124 13555 3196
rect 13485 1036 13555 1124
rect 11220 -1124 11290 -1036
rect 8955 -3284 9025 -3196
rect 6690 -5444 6760 -5356
rect 4425 -7560 4495 -7516
rect 5580 -7560 5650 -7465
rect 6690 -7516 6700 -5444
rect 6750 -7516 6760 -5444
rect 7845 -5495 7915 -5305
rect 8955 -5356 8965 -3284
rect 9015 -5356 9025 -3284
rect 10110 -3335 10180 -3145
rect 11220 -3196 11230 -1124
rect 11280 -3196 11290 -1124
rect 12375 -1175 12445 -985
rect 13485 -1036 13495 1036
rect 13545 -1036 13555 1036
rect 13485 -1124 13555 -1036
rect 11220 -3284 11290 -3196
rect 8955 -5444 9025 -5356
rect 6690 -7560 6760 -7516
rect 7845 -7560 7915 -7465
rect 8955 -7516 8965 -5444
rect 9015 -7516 9025 -5444
rect 10110 -5495 10180 -5305
rect 11220 -5356 11230 -3284
rect 11280 -5356 11290 -3284
rect 12375 -3335 12445 -3145
rect 13485 -3196 13495 -1124
rect 13545 -3196 13555 -1124
rect 13485 -3284 13555 -3196
rect 11220 -5444 11290 -5356
rect 8955 -7560 9025 -7516
rect 10110 -7560 10180 -7465
rect 11220 -7516 11230 -5444
rect 11280 -7516 11290 -5444
rect 12375 -5495 12445 -5305
rect 13485 -5356 13495 -3284
rect 13545 -5356 13555 -3284
rect 13485 -5444 13555 -5356
rect 11220 -7560 11290 -7516
rect 12375 -7560 12445 -7465
rect 13485 -7516 13495 -5444
rect 13545 -7516 13555 -5444
rect 13485 -7560 13555 -7516
<< properties >>
string parameters w 20.00 l 20.00 val 413.6 carea 1.00 cperi 0.17 nx 12 ny 7 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
