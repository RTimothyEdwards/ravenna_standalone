magic
tech EFXH018D
timestamp 1494891594
<< metal2 >>
tri 104 800 264 960 se
tri 264 800 424 960 sw
tri 0 688 104 800 se
rect 104 760 424 800
rect 0 424 104 688
tri 104 640 224 760 nw
tri 304 640 424 760 ne
tri 424 688 528 800 sw
rect 424 424 528 688
rect 0 320 528 424
rect 0 0 104 320
rect 424 0 528 320
<< end >>
