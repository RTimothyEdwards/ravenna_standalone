magic
tech EFXH018D
magscale 1 2
timestamp 1555546584
<< metal2 >>
tri 9 1739 217 1947 se
rect 217 1739 857 1947
tri 857 1739 1065 1947 sw
rect 9 1723 1065 1739
rect 9 1045 217 1723
tri 217 1611 329 1723 nw
tri 745 1611 857 1723 ne
tri 217 1045 329 1157 sw
tri 745 1045 857 1157 se
rect 857 1045 1065 1723
tri 9 838 216 1045 ne
rect 216 838 1065 1045
rect 349 837 697 838
rect 9 235 217 444
tri 217 235 329 347 sw
tri 745 235 857 347 se
rect 857 235 1065 838
tri 9 27 217 235 ne
rect 217 27 857 235
tri 857 27 1065 235 nw
<< end >>
