magic
tech EFXH018D
timestamp 1523029302
<< metal2 >>
tri 0 856 104 960 se
rect 104 856 424 960
tri 424 856 528 960 sw
rect 0 848 528 856
rect 0 496 104 848
tri 104 792 160 848 nw
tri 368 792 424 848 ne
tri 264 576 424 736 se
rect 424 576 528 848
tri 184 496 264 576 se
rect 264 528 528 576
rect 0 416 264 496
tri 264 416 368 528 nw
rect 0 104 104 416
tri 104 256 264 416 nw
tri 104 104 160 160 sw
tri 368 104 424 160 se
rect 424 104 528 528
tri 0 0 104 104 ne
rect 104 0 424 104
tri 424 0 528 104 nw
<< end >>
