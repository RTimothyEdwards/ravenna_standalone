magic
tech EFXH018A
magscale 1 2
timestamp 1527162843
<< checkpaint >>
rect 3694 -2560 10904 4552
<< metal1 >>
rect 5694 2530 5894 2552
rect 5694 2424 8572 2530
rect 5694 2352 5894 2424
rect 6082 2266 6128 2424
rect 6772 2266 6818 2424
rect 7260 2266 7306 2424
rect 7748 2266 7794 2424
rect 8424 2266 8572 2424
rect 6082 1838 6130 2266
rect 6226 1860 6274 2244
rect 6622 2230 6670 2244
rect 6622 1860 6674 2230
rect 6082 1730 6128 1838
rect 5700 1538 5900 1606
rect 6226 1538 6272 1860
rect 5700 1450 6272 1538
rect 5700 1406 5900 1450
rect 6082 850 6130 1278
rect 6226 1256 6272 1450
rect 6628 1256 6674 1860
rect 6766 1838 6818 2266
rect 7108 1860 7156 2244
rect 6772 1726 6818 1838
rect 6226 872 6274 1256
rect 6622 1094 6674 1256
rect 6766 1094 6814 1278
rect 7110 1622 7156 1860
rect 7252 1838 7306 2266
rect 7260 1726 7306 1838
rect 7396 1860 7444 2244
rect 7396 1622 7442 1860
rect 7110 1422 7442 1622
rect 7110 1256 7156 1422
rect 6622 978 6814 1094
rect 6622 872 6674 978
rect 6628 864 6674 872
rect 6766 850 6814 978
rect 7108 872 7156 1256
rect 7252 850 7300 1278
rect 7396 1256 7442 1422
rect 7738 1838 7794 2266
rect 7882 2234 7930 2244
rect 7882 1860 7932 2234
rect 7748 1728 7794 1838
rect 7396 872 7444 1256
rect 7738 1122 7786 1278
rect 7886 1256 7932 1860
rect 8278 1860 8326 2244
rect 7882 1122 7932 1256
rect 7738 1024 7932 1122
rect 7396 868 7442 872
rect 7738 850 7786 1024
rect 7882 872 7932 1024
rect 8278 1412 8324 1860
rect 8422 1838 8572 2266
rect 8424 1490 8572 1838
rect 8698 1720 8864 1808
rect 8698 1520 8898 1720
rect 8704 1412 8904 1422
rect 8278 1324 8904 1412
rect 8278 1256 8324 1324
rect 8278 872 8326 1256
rect 7886 870 7932 872
rect 8278 868 8324 872
rect 8422 850 8470 1278
rect 8704 1222 8904 1324
rect 5702 694 5902 742
rect 6082 694 6128 850
rect 6768 694 6814 850
rect 7254 694 7300 850
rect 7740 694 7786 850
rect 8424 694 8470 850
rect 5702 590 8470 694
rect 5702 588 6222 590
rect 5702 542 5902 588
rect 6006 544 6222 588
rect 8096 588 8470 590
rect 8096 544 8328 588
rect 6006 384 8328 544
rect 6314 248 6378 384
rect 6632 264 6718 384
rect 5702 106 5902 190
rect 5702 28 6068 106
rect 5702 -10 5902 28
rect 6220 24 6354 110
rect 6250 -4 6354 24
rect 6250 -60 6444 -4
rect 6380 -140 6444 -60
rect 7016 226 7086 384
rect 7396 256 7466 384
rect 7776 208 7840 384
rect 5698 -184 5898 -140
rect 6122 -184 6334 -182
rect 5698 -232 6334 -184
rect 6380 -186 6690 -140
rect 5698 -306 6584 -232
rect 6644 -234 6690 -186
rect 6644 -280 6740 -234
rect 5698 -340 5898 -306
rect 7018 -352 7084 -234
rect 7392 -352 7472 -252
rect 7772 -352 7838 -144
rect 8474 -352 8618 540
rect 6088 -512 8618 -352
<< obsm1 >>
rect 6314 2358 6386 2376
rect 6512 2360 6584 2376
rect 6290 2292 6420 2358
rect 6484 2292 6614 2360
rect 6998 2358 7070 2376
rect 6974 2292 7104 2358
rect 7484 2360 7556 2376
rect 7456 2292 7584 2360
rect 7970 2358 8042 2376
rect 8168 2360 8240 2376
rect 7946 2292 8076 2358
rect 8148 2292 8276 2360
rect 6424 1860 6472 2244
rect 6424 1548 6470 1860
rect 6332 1452 6580 1548
rect 6424 1256 6470 1452
rect 6910 2232 6958 2244
rect 6910 1860 7002 2232
rect 6956 1546 7002 1860
rect 6844 1446 7002 1546
rect 6424 872 6472 1256
rect 6956 1256 7002 1446
rect 7594 1860 7642 2244
rect 6910 876 7002 1256
rect 6910 872 6958 876
rect 7594 1546 7640 1860
rect 7594 1446 7740 1546
rect 7594 1256 7640 1446
rect 7594 872 7642 1256
rect 8080 1860 8128 2244
rect 8080 1548 8126 1860
rect 7978 1456 8224 1548
rect 8080 1256 8126 1456
rect 8080 872 8128 1256
rect 6282 744 6416 810
rect 6482 744 6614 810
rect 6314 740 6386 744
rect 6512 740 6584 744
rect 6970 744 7104 810
rect 6998 740 7070 744
rect 7454 744 7586 810
rect 7484 740 7556 744
rect 7942 744 8076 810
rect 8142 744 8304 810
rect 7970 740 8042 744
rect 8168 740 8240 744
rect 6120 202 6196 320
rect 6502 214 6570 326
rect 6120 156 6452 202
rect 6502 168 6782 214
rect 6124 -22 6172 156
rect 6406 122 6452 156
rect 6406 56 6688 122
rect 6124 -136 6200 -22
rect 6736 -22 6782 168
rect 6490 -94 6782 -22
rect 6834 168 6894 326
rect 7204 210 7274 328
rect 7586 252 7652 328
rect 7204 180 7506 210
rect 6834 -34 6888 168
rect 6946 164 7506 180
rect 7586 178 7728 252
rect 7916 322 7974 384
rect 8096 220 8172 334
rect 8234 322 8292 384
rect 6946 134 7250 164
rect 6946 -4 7012 134
rect 6736 -142 6782 -94
rect 6828 -50 6888 -34
rect 7086 -50 7152 88
rect 6828 -96 7152 -50
rect 7200 -46 7250 134
rect 7296 32 7366 118
rect 7448 110 7506 164
rect 7664 110 7728 178
rect 8070 162 8188 220
rect 7434 36 7610 110
rect 7200 -96 7272 -46
rect 7320 -142 7366 32
rect 7664 34 8076 110
rect 7664 -10 7728 34
rect 6736 -188 7366 -142
rect 7582 -92 7728 -10
rect 8132 -25 8188 162
rect 8072 -87 8188 -25
rect 7582 -204 7648 -92
rect 7918 -352 7977 -236
rect 8234 -352 8292 -236
<< metal2 >>
rect 7276 1722 8874 1798
rect 7276 1598 7350 1722
rect 7196 1442 7350 1598
rect 8346 1490 8572 1640
rect 8346 1144 8498 1490
rect 8346 992 8618 1144
rect 8474 388 8618 992
rect 5980 32 6336 102
<< obsm2 >>
rect 5966 2424 8044 2480
rect 5980 678 6048 2424
rect 6316 2282 6388 2424
rect 6512 2226 6584 2368
rect 7000 2282 7072 2424
rect 7484 2226 7556 2368
rect 7972 2282 8044 2424
rect 8176 2226 8248 2368
rect 6178 2170 8248 2226
rect 6180 932 6246 2170
rect 6372 1534 6564 1544
rect 6870 1534 6974 1536
rect 6362 1460 6996 1534
rect 6372 1458 6564 1460
rect 6870 1450 6974 1460
rect 7614 1534 7724 1542
rect 8008 1534 8200 1546
rect 7614 1460 8214 1534
rect 7614 1458 7724 1460
rect 8346 932 8412 934
rect 6180 876 8412 932
rect 6312 734 6384 876
rect 6512 678 6584 820
rect 7000 734 7072 876
rect 7484 678 7556 820
rect 7972 734 8044 876
rect 8172 678 8242 820
rect 5980 622 8242 678
rect 8100 234 8166 622
rect 8346 560 8412 876
rect 8244 494 8412 560
rect 8244 104 8310 494
rect 7898 38 8310 104
<< labels >>
rlabel metal1 6226 872 6274 1256 6 AIN1
port 1 nsew
rlabel metal1 6226 1256 6272 1450 6 AIN1
port 1 nsew
rlabel metal1 5700 1406 5900 1450 6 AIN1
port 1 nsew
rlabel metal1 5700 1450 6272 1538 6 AIN1
port 1 nsew
rlabel metal1 6226 1538 6272 1860 6 AIN1
port 1 nsew
rlabel metal1 5700 1538 5900 1606 6 AIN1
port 1 nsew
rlabel metal1 6226 1860 6274 2244 6 AIN1
port 1 nsew
rlabel metal1 8278 868 8324 872 6 AIN2
port 2 nsew
rlabel metal1 8704 1222 8904 1324 6 AIN2
port 2 nsew
rlabel metal1 8278 872 8326 1256 6 AIN2
port 2 nsew
rlabel metal1 8278 1256 8324 1324 6 AIN2
port 2 nsew
rlabel metal1 8278 1324 8904 1412 6 AIN2
port 2 nsew
rlabel metal1 8704 1412 8904 1422 6 AIN2
port 2 nsew
rlabel metal1 8278 1412 8324 1860 6 AIN2
port 2 nsew
rlabel metal1 8278 1860 8326 2244 6 AIN2
port 2 nsew
rlabel metal2 7196 1442 7350 1598 6 AOUT
port 3 nsew
rlabel metal2 7276 1598 7350 1722 6 AOUT
port 3 nsew
rlabel metal2 7276 1722 8874 1798 6 AOUT
port 3 nsew
rlabel metal1 7396 868 7442 872 6 AOUT
port 3 nsew
rlabel metal1 7396 872 7444 1256 6 AOUT
port 3 nsew
rlabel metal1 7396 1256 7442 1422 6 AOUT
port 3 nsew
rlabel metal1 7108 872 7156 1256 6 AOUT
port 3 nsew
rlabel metal1 7110 1256 7156 1422 6 AOUT
port 3 nsew
rlabel metal1 8698 1520 8898 1720 6 AOUT
port 3 nsew
rlabel metal1 8698 1720 8864 1808 6 AOUT
port 3 nsew
rlabel metal1 7110 1422 7442 1622 6 AOUT
port 3 nsew
rlabel metal1 7396 1622 7442 1860 6 AOUT
port 3 nsew
rlabel metal1 7396 1860 7444 2244 6 AOUT
port 3 nsew
rlabel metal1 7110 1622 7156 1860 6 AOUT
port 3 nsew
rlabel metal1 7108 1860 7156 2244 6 AOUT
port 3 nsew
rlabel metal2 5980 32 6336 102 6 SEL
port 4 nsew
rlabel metal1 6644 -280 6740 -234 8 SEL
port 4 nsew
rlabel metal1 6644 -234 6690 -186 8 SEL
port 4 nsew
rlabel metal1 6380 -186 6690 -140 8 SEL
port 4 nsew
rlabel metal1 6380 -140 6444 -60 8 SEL
port 4 nsew
rlabel metal1 6250 -60 6444 -4 8 SEL
port 4 nsew
rlabel metal1 6250 -4 6354 24 6 SEL
port 4 nsew
rlabel metal1 6220 24 6354 110 6 SEL
port 4 nsew
rlabel metal1 5702 -10 5902 28 6 SEL
port 4 nsew
rlabel metal1 5702 28 6068 106 6 SEL
port 4 nsew
rlabel metal1 5702 106 5902 190 6 SEL
port 4 nsew
rlabel metal1 5698 -340 5898 -306 8 VDD1V8
port 5 nsew
rlabel metal1 5698 -306 6584 -232 8 VDD1V8
port 5 nsew
rlabel metal1 5698 -232 6334 -184 8 VDD1V8
port 5 nsew
rlabel metal1 6122 -184 6334 -182 8 VDD1V8
port 5 nsew
rlabel metal1 5698 -184 5898 -140 8 VDD1V8
port 5 nsew
rlabel metal2 8474 388 8618 992 6 VDD3V3
port 6 nsew
rlabel metal2 8346 992 8618 1144 6 VDD3V3
port 6 nsew
rlabel metal2 8346 1144 8498 1490 6 VDD3V3
port 6 nsew
rlabel metal2 8346 1490 8572 1640 6 VDD3V3
port 6 nsew
rlabel metal1 6088 -512 8618 -352 8 VDD3V3
port 6 nsew
rlabel metal1 8474 -352 8618 540 6 VDD3V3
port 6 nsew
rlabel metal1 7772 -352 7838 -144 8 VDD3V3
port 6 nsew
rlabel metal1 7392 -352 7472 -252 8 VDD3V3
port 6 nsew
rlabel metal1 7018 -352 7084 -234 8 VDD3V3
port 6 nsew
rlabel metal1 8424 1490 8572 1838 6 VDD3V3
port 6 nsew
rlabel metal1 7748 1728 7794 1838 6 VDD3V3
port 6 nsew
rlabel metal1 7260 1726 7306 1838 6 VDD3V3
port 6 nsew
rlabel metal1 6772 1726 6818 1838 6 VDD3V3
port 6 nsew
rlabel metal1 6082 1730 6128 1838 6 VDD3V3
port 6 nsew
rlabel metal1 8422 1838 8572 2266 6 VDD3V3
port 6 nsew
rlabel metal1 7738 1838 7794 2266 6 VDD3V3
port 6 nsew
rlabel metal1 7252 1838 7306 2266 6 VDD3V3
port 6 nsew
rlabel metal1 6766 1838 6818 2266 6 VDD3V3
port 6 nsew
rlabel metal1 6082 1838 6130 2266 6 VDD3V3
port 6 nsew
rlabel metal1 8424 2266 8572 2424 6 VDD3V3
port 6 nsew
rlabel metal1 7748 2266 7794 2424 6 VDD3V3
port 6 nsew
rlabel metal1 7260 2266 7306 2424 6 VDD3V3
port 6 nsew
rlabel metal1 6772 2266 6818 2424 6 VDD3V3
port 6 nsew
rlabel metal1 6082 2266 6128 2424 6 VDD3V3
port 6 nsew
rlabel metal1 5694 2352 5894 2424 6 VDD3V3
port 6 nsew
rlabel metal1 5694 2424 8572 2530 6 VDD3V3
port 6 nsew
rlabel metal1 5694 2530 5894 2552 6 VDD3V3
port 6 nsew
rlabel metal1 7776 208 7840 384 6 VSSA
port 7 nsew
rlabel metal1 7396 256 7466 384 6 VSSA
port 7 nsew
rlabel metal1 7016 226 7086 384 6 VSSA
port 7 nsew
rlabel metal1 6632 264 6718 384 6 VSSA
port 7 nsew
rlabel metal1 6314 248 6378 384 6 VSSA
port 7 nsew
rlabel metal1 6006 384 8328 544 6 VSSA
port 7 nsew
rlabel metal1 8096 544 8328 588 6 VSSA
port 7 nsew
rlabel metal1 8096 588 8470 590 6 VSSA
port 7 nsew
rlabel metal1 6006 544 6222 588 6 VSSA
port 7 nsew
rlabel metal1 5702 542 5902 588 6 VSSA
port 7 nsew
rlabel metal1 5702 588 6222 590 6 VSSA
port 7 nsew
rlabel metal1 5702 590 8470 694 6 VSSA
port 7 nsew
rlabel metal1 8424 694 8470 850 6 VSSA
port 7 nsew
rlabel metal1 7740 694 7786 850 6 VSSA
port 7 nsew
rlabel metal1 7254 694 7300 850 6 VSSA
port 7 nsew
rlabel metal1 6768 694 6814 850 6 VSSA
port 7 nsew
rlabel metal1 6082 694 6128 850 6 VSSA
port 7 nsew
rlabel metal1 5702 694 5902 742 6 VSSA
port 7 nsew
rlabel metal1 8422 850 8470 1278 6 VSSA
port 7 nsew
rlabel metal1 7886 870 7932 872 6 VSSA
port 7 nsew
rlabel metal1 7882 872 7932 1024 6 VSSA
port 7 nsew
rlabel metal1 7738 850 7786 1024 6 VSSA
port 7 nsew
rlabel metal1 7738 1024 7932 1122 6 VSSA
port 7 nsew
rlabel metal1 7882 1122 7932 1256 6 VSSA
port 7 nsew
rlabel metal1 7886 1256 7932 1860 6 VSSA
port 7 nsew
rlabel metal1 7738 1122 7786 1278 6 VSSA
port 7 nsew
rlabel metal1 7252 850 7300 1278 6 VSSA
port 7 nsew
rlabel metal1 6766 850 6814 978 6 VSSA
port 7 nsew
rlabel metal1 6628 864 6674 872 6 VSSA
port 7 nsew
rlabel metal1 6622 872 6674 978 6 VSSA
port 7 nsew
rlabel metal1 6622 978 6814 1094 6 VSSA
port 7 nsew
rlabel metal1 6766 1094 6814 1278 6 VSSA
port 7 nsew
rlabel metal1 6622 1094 6674 1256 6 VSSA
port 7 nsew
rlabel metal1 6628 1256 6674 1860 6 VSSA
port 7 nsew
rlabel metal1 6082 850 6130 1278 6 VSSA
port 7 nsew
rlabel metal1 7882 1860 7932 2234 6 VSSA
port 7 nsew
rlabel metal1 6622 1860 6674 2230 6 VSSA
port 7 nsew
rlabel metal1 7882 2234 7930 2244 6 VSSA
port 7 nsew
rlabel metal1 6622 2230 6670 2244 6 VSSA
port 7 nsew
<< properties >>
string LEFview TRUE
string FIXED_BBOX 5694 -560 8904 2552
string GDS_FILE ~/design/ip/AMUX2_3V/10.0/gds/AMUX2_3V.gds
string GDS_START 24452
string GDS_END 35244
<< end >>
