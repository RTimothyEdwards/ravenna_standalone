magic
tech EFXH018D
timestamp 1494891594
<< metal2 >>
tri 16 848 128 960 se
rect 128 864 424 960
tri 424 864 528 960 sw
rect 128 848 528 864
rect 16 608 128 848
tri 128 800 176 848 nw
tri 368 800 416 848 ne
rect 416 768 528 848
tri 16 496 128 608 ne
tri 128 544 240 656 sw
rect 128 496 416 544
tri 128 432 192 496 ne
rect 192 432 416 496
tri 416 432 528 544 sw
tri 368 384 416 432 ne
rect 16 112 128 208
tri 128 112 176 160 sw
tri 368 112 416 160 se
rect 416 112 528 432
tri 16 0 128 112 ne
rect 128 0 416 112
tri 416 0 528 112 nw
<< end >>
