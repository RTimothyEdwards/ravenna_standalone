magic
tech EFXH018D
magscale 1 2
timestamp 1567005482
<< metal1 >>
rect 16408 20636 16460 20692
rect 16516 20636 16616 20692
rect 16672 20636 16772 20692
rect 16828 20636 16928 20692
rect 16984 20636 17084 20692
rect 17140 20636 17192 20692
rect 4106 20468 4116 20524
rect 4172 20468 4182 20524
rect 4106 20422 4182 20468
rect 3322 20356 3332 20412
rect 3388 20356 3398 20412
rect 20458 20356 20468 20412
rect 20524 20356 20534 20412
rect 2538 20244 2548 20300
rect 2604 20244 2614 20300
rect 3658 20244 3668 20300
rect 3724 20244 3734 20300
rect 3994 20264 4004 20320
rect 4060 20264 4070 20320
rect 4452 20300 4508 20310
rect 5012 20300 5068 20310
rect 4330 20244 4340 20300
rect 4396 20244 4406 20300
rect 4666 20244 4676 20300
rect 4732 20244 4742 20300
rect 4452 20234 4508 20244
rect 5012 20234 5068 20244
rect 5348 20300 5404 20310
rect 11956 20300 12012 20310
rect 14084 20300 14140 20310
rect 6010 20244 6020 20300
rect 6076 20244 6086 20300
rect 6346 20244 6356 20300
rect 6412 20244 6422 20300
rect 10266 20244 10276 20300
rect 10332 20244 10342 20300
rect 12282 20244 12292 20300
rect 12348 20244 12358 20300
rect 5348 20234 5404 20244
rect 11956 20234 12012 20244
rect 14084 20234 14140 20244
rect 14308 20300 14364 20310
rect 19348 20300 19404 20310
rect 18106 20244 18116 20300
rect 18172 20244 18182 20300
rect 14308 20234 14364 20244
rect 19348 20234 19404 20244
rect 21140 20300 21196 20310
rect 21140 20234 21196 20244
rect 22372 20300 22428 20310
rect 22372 20234 22428 20244
rect 23156 20300 23212 20310
rect 23156 20234 23212 20244
rect 3780 20188 3836 20198
rect 12740 20188 12796 20198
rect 1082 20132 1092 20188
rect 1148 20132 1158 20188
rect 1306 20132 1316 20188
rect 1372 20132 1382 20188
rect 4106 20132 4116 20188
rect 4172 20132 4182 20188
rect 8810 20132 8820 20188
rect 8876 20132 8886 20188
rect 9034 20132 9044 20188
rect 9100 20132 9110 20188
rect 10938 20132 10948 20188
rect 11004 20132 11014 20188
rect 3780 20122 3836 20132
rect 4900 20076 4966 20126
rect 12740 20122 12796 20132
rect 13076 20188 13132 20198
rect 13626 20132 13636 20188
rect 13692 20132 13702 20188
rect 16762 20132 16772 20188
rect 16828 20132 16838 20188
rect 16986 20132 16996 20188
rect 17052 20132 17062 20188
rect 18778 20132 18788 20188
rect 18844 20132 18854 20188
rect 19898 20183 19908 20188
rect 19801 20137 19908 20183
rect 19898 20132 19908 20137
rect 19964 20132 19974 20188
rect 13076 20122 13132 20132
rect 4890 20020 4900 20076
rect 4956 20020 4966 20076
rect 6234 20076 6310 20117
rect 6234 20020 6244 20076
rect 6300 20020 6310 20076
rect 21466 20076 21542 20163
rect 22250 20132 22260 20188
rect 22316 20132 22326 20188
rect 21466 20020 21476 20076
rect 21532 20020 21542 20076
rect 22810 20076 22886 20117
rect 22810 20020 22820 20076
rect 22876 20020 22886 20076
rect 23482 20076 23558 20117
rect 23482 20020 23492 20076
rect 23548 20020 23558 20076
rect 13300 19964 13356 19974
rect 12842 19908 12852 19964
rect 12908 19908 12918 19964
rect 13300 19898 13356 19908
rect 5992 19740 6044 19796
rect 6100 19740 6200 19796
rect 6256 19740 6356 19796
rect 6412 19740 6512 19796
rect 6568 19740 6668 19796
rect 6724 19740 6776 19796
rect 4228 19628 4284 19638
rect 21578 19623 21588 19628
rect 4228 19562 4284 19572
rect 21466 19572 21588 19623
rect 21644 19572 21654 19628
rect 21466 19524 21542 19572
rect 22698 19552 22820 19608
rect 22876 19552 22886 19608
rect 22698 19524 22774 19552
rect 19338 19460 19348 19516
rect 19404 19460 19414 19516
rect 19338 19423 19414 19460
rect 1988 19404 2044 19414
rect 12628 19404 12684 19414
rect 1866 19348 1876 19404
rect 1932 19348 1942 19404
rect 2986 19348 2996 19404
rect 3052 19348 3062 19404
rect 9146 19348 9156 19404
rect 9212 19348 9222 19404
rect 9370 19348 9380 19404
rect 9436 19348 9446 19404
rect 11610 19348 11620 19404
rect 11676 19348 11686 19404
rect 1988 19338 2044 19348
rect 12628 19338 12684 19348
rect 12740 19404 12796 19414
rect 15418 19348 15428 19404
rect 15484 19348 15494 19404
rect 15642 19348 15652 19404
rect 15708 19348 15718 19404
rect 12740 19338 12796 19348
rect 4116 19292 4172 19302
rect 4564 19292 4620 19302
rect 4172 19241 4279 19287
rect 4442 19236 4452 19292
rect 4508 19236 4518 19292
rect 4778 19256 4788 19312
rect 4844 19256 4854 19312
rect 19124 19292 19180 19302
rect 19796 19292 19852 19302
rect 5129 19264 5287 19287
rect 4116 19226 4172 19236
rect 4564 19226 4620 19236
rect 5114 19241 5287 19264
rect 84 19180 140 19190
rect 5114 19180 5190 19241
rect 5338 19236 5348 19292
rect 5404 19236 5414 19292
rect 8026 19236 8036 19292
rect 8092 19236 8102 19292
rect 16762 19236 16772 19292
rect 16828 19236 16838 19292
rect 18778 19236 18788 19292
rect 18844 19236 18854 19292
rect 19450 19236 19460 19292
rect 19516 19236 19526 19292
rect 21588 19292 21644 19302
rect 20025 19241 20183 19287
rect 19124 19226 19180 19236
rect 19796 19226 19852 19236
rect 21588 19226 21644 19236
rect 22820 19292 22876 19302
rect 22820 19226 22876 19236
rect 11060 19180 11116 19190
rect 20692 19180 20748 19190
rect 3882 19124 3892 19180
rect 3948 19124 3958 19180
rect 5114 19124 5124 19180
rect 5180 19124 5190 19180
rect 7130 19124 7140 19180
rect 7196 19124 7206 19180
rect 17434 19124 17444 19180
rect 17500 19124 17510 19180
rect 20585 19129 20692 19175
rect 84 19114 140 19124
rect 4778 19068 4854 19124
rect 11060 19114 11116 19124
rect 20692 19114 20748 19124
rect 20804 19180 20860 19190
rect 22148 19180 22204 19190
rect 22041 19129 22148 19175
rect 20804 19114 20860 19124
rect 23594 19175 23604 19180
rect 23273 19129 23604 19175
rect 23594 19124 23604 19129
rect 23660 19124 23670 19180
rect 22148 19114 22204 19124
rect 4778 19012 4788 19068
rect 4844 19012 4854 19068
rect 16408 18844 16460 18900
rect 16516 18844 16616 18900
rect 16672 18844 16772 18900
rect 16828 18844 16928 18900
rect 16984 18844 17084 18900
rect 17140 18844 17192 18900
rect 410 18676 420 18732
rect 476 18676 486 18732
rect 4106 18676 4116 18732
rect 4172 18676 4182 18732
rect 74 18569 84 18625
rect 140 18569 150 18625
rect 4106 18620 4182 18676
rect 4890 18676 4900 18732
rect 4956 18676 4966 18732
rect 4890 18630 4966 18676
rect 7354 18676 7364 18732
rect 7420 18676 7430 18732
rect 7354 18630 7430 18676
rect 11834 18676 11844 18732
rect 11900 18676 11910 18732
rect 5796 18620 5852 18630
rect 74 18486 150 18569
rect 11834 18582 11910 18676
rect 12394 18676 12404 18732
rect 12460 18676 12470 18732
rect 12394 18582 12470 18676
rect 15306 18676 15316 18732
rect 15372 18676 15382 18732
rect 15306 18630 15382 18676
rect 20346 18615 20356 18620
rect 20249 18569 20356 18615
rect 20346 18564 20356 18569
rect 20412 18564 20422 18620
rect 21690 18615 21700 18620
rect 21593 18569 21700 18615
rect 21690 18564 21700 18569
rect 21756 18564 21766 18620
rect 5796 18554 5852 18564
rect 1988 18508 2044 18518
rect 3780 18508 3836 18518
rect 746 18452 756 18508
rect 812 18452 822 18508
rect 2650 18452 2660 18508
rect 2716 18452 2772 18508
rect 3434 18452 3444 18508
rect 3500 18452 3510 18508
rect 3612 18452 3668 18508
rect 3724 18452 3734 18508
rect 4452 18508 4508 18518
rect 5124 18508 5180 18518
rect 5572 18508 5628 18518
rect 6244 18508 6300 18518
rect 4121 18457 4279 18503
rect 1988 18442 2044 18452
rect 3780 18442 3836 18452
rect 4666 18452 4676 18508
rect 4732 18452 4742 18508
rect 5226 18452 5236 18508
rect 5292 18452 5302 18508
rect 5674 18452 5684 18508
rect 5740 18452 5750 18508
rect 6122 18452 6132 18508
rect 6188 18452 6198 18508
rect 4452 18442 4508 18452
rect 5124 18442 5180 18452
rect 5572 18442 5628 18452
rect 6244 18442 6300 18452
rect 6356 18508 6412 18518
rect 6356 18442 6412 18452
rect 6468 18508 6524 18518
rect 6468 18442 6524 18452
rect 7588 18508 7644 18518
rect 11620 18508 11676 18518
rect 7690 18452 7700 18508
rect 7756 18452 7766 18508
rect 10266 18452 10276 18508
rect 10332 18452 10342 18508
rect 7588 18442 7644 18452
rect 11620 18442 11676 18452
rect 12740 18508 12796 18518
rect 19796 18508 19852 18518
rect 13417 18457 13575 18503
rect 14522 18452 14532 18508
rect 14588 18452 14598 18508
rect 14746 18452 14756 18508
rect 14812 18452 14822 18508
rect 15046 18452 15092 18508
rect 15148 18452 15158 18508
rect 17322 18452 17332 18508
rect 17388 18452 17398 18508
rect 12740 18442 12796 18452
rect 3108 18396 3164 18406
rect 13748 18396 13814 18446
rect 19796 18442 19852 18452
rect 20468 18508 20524 18518
rect 20468 18442 20524 18452
rect 21140 18508 21196 18518
rect 21140 18442 21196 18452
rect 21812 18508 21868 18518
rect 21812 18442 21868 18452
rect 22484 18508 22540 18518
rect 22484 18442 22540 18452
rect 4890 18340 4900 18396
rect 4956 18340 4966 18396
rect 5898 18340 5908 18396
rect 5964 18340 5974 18396
rect 7354 18340 7364 18396
rect 7420 18340 7430 18396
rect 8922 18340 8932 18396
rect 8988 18340 8998 18396
rect 9146 18340 9156 18396
rect 9212 18340 9222 18396
rect 10938 18340 10948 18396
rect 11004 18340 11014 18396
rect 13738 18340 13748 18396
rect 13804 18340 13814 18396
rect 14410 18340 14420 18396
rect 14476 18340 14486 18396
rect 16538 18340 16548 18396
rect 16604 18340 16614 18396
rect 18442 18340 18452 18396
rect 18508 18340 18518 18396
rect 18666 18340 18676 18396
rect 18732 18340 18742 18396
rect 23146 18340 23156 18396
rect 23212 18340 23222 18396
rect 3108 18330 3164 18340
rect 1530 18284 1606 18325
rect 186 18228 196 18284
rect 252 18228 262 18284
rect 1530 18228 1540 18284
rect 1596 18228 1606 18284
rect 4106 18284 4182 18334
rect 4106 18228 4116 18284
rect 4172 18228 4182 18284
rect 4554 18284 4630 18325
rect 4554 18228 4564 18284
rect 4620 18228 4630 18284
rect 12282 18284 12358 18325
rect 12282 18228 12292 18284
rect 12348 18228 12358 18284
rect 12954 18284 13030 18325
rect 12954 18228 12964 18284
rect 13020 18228 13030 18284
rect 20906 18284 20982 18325
rect 20906 18228 20916 18284
rect 20972 18228 20982 18284
rect 22250 18284 22326 18325
rect 22250 18228 22260 18284
rect 22316 18228 22326 18284
rect 22922 18284 22998 18325
rect 22922 18228 22932 18284
rect 22988 18228 22998 18284
rect 5992 17948 6044 18004
rect 6100 17948 6200 18004
rect 6256 17948 6356 18004
rect 6412 17948 6512 18004
rect 6568 17948 6668 18004
rect 6724 17948 6776 18004
rect 19002 17668 19012 17724
rect 19068 17668 19078 17724
rect 19002 17627 19078 17668
rect 4228 17612 4284 17622
rect 6794 17556 6804 17612
rect 6860 17556 6870 17612
rect 7018 17556 7028 17612
rect 7084 17556 7094 17612
rect 11050 17556 11060 17612
rect 11116 17556 11126 17612
rect 11274 17556 11284 17612
rect 11340 17556 11350 17612
rect 15418 17556 15428 17612
rect 15484 17556 15494 17612
rect 15642 17556 15652 17612
rect 15708 17556 15718 17612
rect 4228 17546 4284 17556
rect 420 17500 476 17510
rect 2548 17500 2604 17510
rect 1642 17444 1652 17500
rect 1708 17444 1718 17500
rect 2090 17444 2100 17500
rect 2156 17444 2166 17500
rect 420 17434 476 17444
rect 2548 17434 2604 17444
rect 2660 17500 2716 17510
rect 3220 17500 3276 17510
rect 3668 17500 3724 17510
rect 20244 17500 20300 17510
rect 2716 17449 2823 17495
rect 3098 17444 3108 17500
rect 3164 17444 3174 17500
rect 3546 17444 3556 17500
rect 3612 17444 3622 17500
rect 4106 17444 4116 17500
rect 4172 17444 4182 17500
rect 8250 17444 8260 17500
rect 8316 17444 8326 17500
rect 9370 17444 9380 17500
rect 9436 17444 9446 17500
rect 9670 17444 9716 17500
rect 9772 17444 9782 17500
rect 12394 17444 12404 17500
rect 12460 17444 12470 17500
rect 16874 17444 16884 17500
rect 16940 17444 16950 17500
rect 2660 17434 2716 17444
rect 3220 17434 3276 17444
rect 3668 17434 3724 17444
rect 20244 17434 20300 17444
rect 21476 17500 21532 17510
rect 21476 17434 21532 17444
rect 22708 17500 22764 17510
rect 22708 17434 22764 17444
rect 196 17388 252 17398
rect 9940 17388 9996 17398
rect 18778 17388 18854 17434
rect 20804 17388 20860 17398
rect 9034 17332 9044 17388
rect 9100 17332 9110 17388
rect 13290 17332 13300 17388
rect 13356 17332 13366 17388
rect 17658 17332 17668 17388
rect 17724 17332 17734 17388
rect 18778 17332 18788 17388
rect 18844 17332 18854 17388
rect 19562 17332 19572 17388
rect 19628 17332 19638 17388
rect 20697 17337 20804 17383
rect 21354 17332 21364 17388
rect 21420 17332 21430 17388
rect 22026 17383 22036 17388
rect 21929 17337 22036 17383
rect 22026 17332 22036 17337
rect 22092 17332 22102 17388
rect 22586 17332 22596 17388
rect 22652 17332 22662 17388
rect 23706 17383 23716 17388
rect 23161 17337 23716 17383
rect 23706 17332 23716 17337
rect 23772 17332 23782 17388
rect 196 17322 252 17332
rect 746 17266 822 17323
rect 1876 17276 1942 17326
rect 746 17210 756 17266
rect 812 17210 822 17266
rect 1866 17220 1876 17276
rect 1932 17220 1942 17276
rect 2314 17276 2390 17322
rect 2314 17220 2324 17276
rect 2380 17220 2390 17276
rect 3098 17276 3174 17332
rect 3098 17220 3108 17276
rect 3164 17220 3174 17276
rect 3220 17276 3296 17332
rect 3892 17276 3958 17326
rect 9940 17322 9996 17332
rect 20804 17322 20860 17332
rect 3220 17225 3230 17276
rect 3286 17225 3296 17276
rect 3882 17220 3892 17276
rect 3948 17220 3958 17276
rect 3230 17210 3286 17220
rect 16408 17052 16460 17108
rect 16516 17052 16616 17108
rect 16672 17052 16772 17108
rect 16828 17052 16928 17108
rect 16984 17052 17084 17108
rect 17140 17052 17192 17108
rect 8810 16884 8820 16940
rect 8876 16884 8886 16940
rect 9482 16884 9492 16940
rect 9548 16884 9558 16940
rect 8810 16837 8886 16884
rect 9492 16834 9558 16884
rect 11050 16884 11060 16940
rect 11116 16884 11126 16940
rect 11050 16838 11126 16884
rect 14746 16884 14756 16940
rect 14812 16884 14822 16940
rect 14746 16838 14822 16884
rect 16874 16884 16884 16940
rect 16940 16884 16950 16940
rect 16874 16838 16950 16884
rect 14644 16828 14700 16838
rect 4192 16772 4228 16828
rect 4284 16772 4294 16828
rect 23370 16772 23380 16828
rect 23436 16772 23446 16828
rect 14644 16762 14700 16772
rect 644 16716 700 16726
rect 644 16650 700 16660
rect 1540 16716 1596 16726
rect 1764 16716 1820 16726
rect 2212 16716 2268 16726
rect 1642 16660 1652 16716
rect 1708 16660 1718 16716
rect 2090 16660 2100 16716
rect 2156 16660 2166 16716
rect 1540 16650 1596 16660
rect 1764 16650 1820 16660
rect 2212 16650 2268 16660
rect 2324 16716 2380 16726
rect 2324 16650 2380 16660
rect 2436 16716 2492 16726
rect 3556 16716 3612 16726
rect 2436 16650 2492 16660
rect 2538 16645 2548 16701
rect 2604 16645 2614 16701
rect 2874 16660 2884 16716
rect 2940 16660 2950 16716
rect 3780 16716 3836 16726
rect 4564 16716 4620 16726
rect 5908 16716 5964 16726
rect 3882 16660 3892 16716
rect 3948 16660 3958 16716
rect 4106 16660 4116 16716
rect 4172 16660 4182 16716
rect 4457 16665 4564 16711
rect 5450 16660 5460 16716
rect 5516 16660 5526 16716
rect 3780 16650 3836 16660
rect 4564 16650 4620 16660
rect 5908 16650 5964 16660
rect 6020 16716 6076 16726
rect 6020 16650 6076 16660
rect 7364 16716 7420 16726
rect 7364 16650 7420 16660
rect 7588 16716 7644 16726
rect 7588 16650 7644 16660
rect 7700 16716 7756 16726
rect 7700 16650 7756 16660
rect 7924 16716 7980 16726
rect 8377 16716 8433 16726
rect 8138 16660 8148 16716
rect 8204 16660 8214 16716
rect 7924 16650 7980 16660
rect 8377 16650 8433 16660
rect 8489 16716 8545 16726
rect 8489 16650 8545 16660
rect 8932 16716 8988 16726
rect 9034 16660 9044 16716
rect 9100 16660 9110 16716
rect 9258 16660 9268 16716
rect 9324 16660 9334 16716
rect 9706 16670 9716 16726
rect 9772 16670 9782 16726
rect 10836 16716 10892 16726
rect 14980 16716 15036 16726
rect 14074 16660 14084 16716
rect 14140 16660 14150 16716
rect 8932 16650 8988 16660
rect 10836 16650 10892 16660
rect 14980 16650 15036 16660
rect 16660 16716 16716 16726
rect 16660 16650 16716 16660
rect 22260 16716 22316 16726
rect 22260 16650 22316 16660
rect 5348 16604 5404 16614
rect 1082 16492 1158 16579
rect 1866 16548 1876 16604
rect 1932 16548 1942 16604
rect 5786 16548 5796 16604
rect 5852 16548 5862 16604
rect 9828 16599 9884 16609
rect 5348 16538 5404 16548
rect 7242 16543 7252 16599
rect 7308 16543 7318 16599
rect 9828 16533 9884 16543
rect 10276 16604 10332 16614
rect 15540 16604 15596 16614
rect 12730 16548 12740 16604
rect 12796 16548 12806 16604
rect 12954 16548 12964 16604
rect 13020 16548 13030 16604
rect 10276 16538 10332 16548
rect 15540 16538 15596 16548
rect 16100 16604 16156 16614
rect 16100 16538 16156 16548
rect 19348 16604 19404 16614
rect 19348 16538 19404 16548
rect 19460 16604 19516 16614
rect 20458 16548 20468 16604
rect 20524 16548 20534 16604
rect 21130 16548 21140 16604
rect 21196 16548 21206 16604
rect 22138 16548 22148 16604
rect 22204 16548 22214 16604
rect 19460 16538 19516 16548
rect 1082 16436 1092 16492
rect 1148 16436 1158 16492
rect 2762 16492 2838 16533
rect 2762 16436 2772 16492
rect 2828 16436 2838 16492
rect 6804 16492 6860 16502
rect 6906 16487 6982 16533
rect 6860 16441 6982 16487
rect 22698 16492 22774 16533
rect 22698 16436 22708 16492
rect 22764 16436 22774 16492
rect 6804 16426 6860 16436
rect 3556 16380 3612 16390
rect 3556 16314 3612 16324
rect 10052 16380 10108 16390
rect 15642 16324 15652 16380
rect 15708 16324 15718 16380
rect 15769 16329 15927 16375
rect 10052 16314 10108 16324
rect 5992 16156 6044 16212
rect 6100 16156 6200 16212
rect 6256 16156 6356 16212
rect 6412 16156 6512 16212
rect 6568 16156 6668 16212
rect 6724 16156 6776 16212
rect 5796 16044 5852 16054
rect 5796 15978 5852 15988
rect 6356 16044 6412 16054
rect 6356 15978 6412 15988
rect 13748 16044 13804 16054
rect 13748 15978 13804 15988
rect 4330 15876 4340 15932
rect 4396 15876 4406 15932
rect 7802 15927 7812 15932
rect 7578 15881 7812 15927
rect 1082 15764 1092 15820
rect 1148 15764 1158 15820
rect 2874 15764 2884 15820
rect 2940 15764 2950 15820
rect 3098 15764 3108 15820
rect 3164 15764 3174 15820
rect 7578 15789 7654 15881
rect 7802 15876 7812 15881
rect 7868 15876 7878 15932
rect 12730 15876 12740 15932
rect 12796 15876 12806 15932
rect 12730 15835 12806 15876
rect 20346 15876 20356 15932
rect 20412 15876 20422 15932
rect 13524 15820 13580 15830
rect 18788 15820 18844 15830
rect 9258 15764 9268 15820
rect 9324 15764 9334 15820
rect 9482 15764 9492 15820
rect 9548 15764 9558 15820
rect 17770 15764 17780 15820
rect 17836 15764 17846 15820
rect 18890 15764 18900 15820
rect 18956 15764 18966 15820
rect 20346 15789 20422 15876
rect 13524 15754 13580 15764
rect 18788 15754 18844 15764
rect 6132 15708 6188 15718
rect 15092 15708 15148 15718
rect 1642 15652 1652 15708
rect 1708 15652 1718 15708
rect 4890 15652 4900 15708
rect 4956 15652 4966 15708
rect 5338 15652 5348 15708
rect 5404 15652 5460 15708
rect 5562 15652 5572 15708
rect 5628 15652 5638 15708
rect 5786 15652 5796 15708
rect 5852 15652 5862 15708
rect 6010 15652 6020 15708
rect 6076 15652 6086 15708
rect 6346 15652 6356 15708
rect 6412 15652 6422 15708
rect 7354 15652 7364 15708
rect 7420 15652 7430 15708
rect 7578 15652 7588 15708
rect 7644 15652 7654 15708
rect 10714 15652 10724 15708
rect 10780 15652 10790 15708
rect 11946 15652 11956 15708
rect 12012 15652 12022 15708
rect 13066 15652 13076 15708
rect 13132 15652 13142 15708
rect 6132 15642 6188 15652
rect 15092 15642 15148 15652
rect 20132 15708 20188 15718
rect 20132 15642 20188 15652
rect 21252 15708 21308 15718
rect 21252 15642 21308 15652
rect 21812 15713 21868 15723
rect 23156 15708 23212 15718
rect 21868 15657 21975 15703
rect 21812 15647 21868 15657
rect 23156 15642 23212 15652
rect 4218 15540 4228 15596
rect 4284 15591 4294 15596
rect 4284 15545 4391 15591
rect 4284 15540 4294 15545
rect 4554 15540 4564 15596
rect 4620 15540 4630 15596
rect 11498 15540 11508 15596
rect 11564 15540 11574 15596
rect 14634 15540 14644 15596
rect 14700 15591 14710 15596
rect 14700 15545 14807 15591
rect 14700 15540 14710 15545
rect 17210 15540 17220 15596
rect 17276 15540 17286 15596
rect 21130 15540 21140 15596
rect 21196 15540 21206 15596
rect 21812 15591 21868 15601
rect 22484 15596 22540 15606
rect 21705 15545 21812 15591
rect 22377 15545 22484 15591
rect 11834 15484 11910 15530
rect 21812 15525 21868 15535
rect 23034 15540 23044 15596
rect 23100 15540 23110 15596
rect 23706 15591 23716 15596
rect 23609 15545 23716 15591
rect 23706 15540 23716 15545
rect 23772 15540 23782 15596
rect 22484 15530 22540 15540
rect 11834 15428 11844 15484
rect 11900 15428 11910 15484
rect 16408 15260 16460 15316
rect 16516 15260 16616 15316
rect 16672 15260 16772 15316
rect 16828 15260 16928 15316
rect 16984 15260 17084 15316
rect 17140 15260 17192 15316
rect 746 15092 756 15148
rect 812 15092 822 15148
rect 1978 15092 1988 15148
rect 2044 15092 2054 15148
rect 4778 15092 4788 15148
rect 4844 15092 4854 15148
rect 756 15045 822 15092
rect 634 15031 644 15036
rect 537 14985 644 15031
rect 634 14980 644 14985
rect 700 14980 710 15036
rect 3642 14980 3668 15036
rect 3724 14980 3734 15036
rect 4345 14995 4452 15051
rect 4508 14995 4518 15051
rect 4778 15046 4854 15092
rect 10378 15092 10388 15148
rect 10444 15092 10454 15148
rect 20122 15092 20132 15148
rect 20188 15092 20198 15148
rect 21690 15092 21700 15148
rect 21756 15092 21766 15148
rect 10378 15054 10454 15092
rect 22932 15041 22988 15051
rect 6458 14980 6468 15036
rect 6524 14980 6534 15036
rect 14298 14980 14308 15036
rect 14364 14980 14374 15036
rect 21130 14980 21140 15036
rect 21196 14980 21206 15036
rect 22825 14985 22932 15031
rect 23604 15036 23660 15046
rect 23497 14985 23604 15031
rect 14298 14934 14374 14980
rect 22932 14975 22988 14985
rect 23604 14970 23660 14980
rect 84 14924 140 14934
rect 84 14858 140 14868
rect 196 14924 252 14934
rect 196 14858 252 14868
rect 1316 14924 1372 14934
rect 1652 14924 1708 14934
rect 2660 14924 2716 14934
rect 1418 14868 1428 14924
rect 1484 14868 1494 14924
rect 2426 14868 2436 14924
rect 2492 14868 2502 14924
rect 1316 14858 1372 14868
rect 1652 14858 1708 14868
rect 2660 14858 2716 14868
rect 3220 14924 3276 14934
rect 4564 14924 4620 14934
rect 22372 14924 22428 14934
rect 4106 14868 4116 14924
rect 4172 14868 4182 14924
rect 7242 14868 7252 14924
rect 7308 14868 7318 14924
rect 9930 14868 9940 14924
rect 9996 14868 10006 14924
rect 11722 14868 11732 14924
rect 11788 14868 11798 14924
rect 18330 14868 18340 14924
rect 18396 14868 18406 14924
rect 3220 14858 3276 14868
rect 4564 14858 4620 14868
rect 22372 14858 22428 14868
rect 22932 14919 22988 14929
rect 22988 14873 23095 14919
rect 22932 14853 22988 14863
rect 10052 14812 10108 14822
rect 1082 14756 1092 14812
rect 1148 14756 1158 14812
rect 2762 14756 2772 14812
rect 2828 14756 2838 14812
rect 4778 14756 4788 14812
rect 4844 14756 4854 14812
rect 3780 14700 3836 14710
rect 3561 14649 3780 14695
rect 6794 14700 6870 14787
rect 8474 14756 8484 14812
rect 8540 14756 8550 14812
rect 8698 14756 8708 14812
rect 8764 14756 8774 14812
rect 10490 14756 10500 14812
rect 10556 14756 10566 14812
rect 12954 14756 12964 14812
rect 13020 14756 13030 14812
rect 13178 14756 13188 14812
rect 13244 14756 13254 14812
rect 16986 14756 16996 14812
rect 17052 14756 17062 14812
rect 17210 14756 17220 14812
rect 17276 14756 17286 14812
rect 19002 14756 19012 14812
rect 19068 14756 19078 14812
rect 10052 14746 10108 14756
rect 6794 14644 6804 14700
rect 6860 14644 6870 14700
rect 11172 14700 11228 14710
rect 14522 14700 14598 14741
rect 11228 14649 11335 14695
rect 14522 14644 14532 14700
rect 14588 14644 14598 14700
rect 3780 14634 3836 14644
rect 11172 14634 11228 14644
rect 5992 14364 6044 14420
rect 6100 14364 6200 14420
rect 6256 14364 6356 14420
rect 6412 14364 6512 14420
rect 6568 14364 6668 14420
rect 6724 14364 6776 14420
rect 9380 14252 9436 14262
rect 4905 14201 5063 14247
rect 9380 14186 9436 14196
rect 3098 14089 3108 14145
rect 3164 14089 3174 14145
rect 3098 14043 3174 14089
rect 4218 14084 4228 14140
rect 4284 14084 4294 14140
rect 6122 14084 6132 14140
rect 6188 14084 6198 14140
rect 6122 14043 6198 14084
rect 8362 14084 8372 14140
rect 8428 14084 8438 14140
rect 8362 14043 8438 14084
rect 16202 14084 16212 14140
rect 16268 14084 16278 14140
rect 16202 14043 16268 14084
rect 3892 14028 3948 14038
rect 5236 14028 5292 14038
rect 18788 14028 18844 14038
rect 1082 13972 1092 14028
rect 1148 13972 1158 14028
rect 1306 13972 1316 14028
rect 1372 13972 1382 14028
rect 3322 13972 3332 14028
rect 3388 13972 3398 14028
rect 4890 13972 4900 14028
rect 4956 13972 4966 14028
rect 7914 13972 7924 14028
rect 7980 13972 7990 14028
rect 12730 13972 12740 14028
rect 12796 13972 12806 14028
rect 3892 13962 3948 13972
rect 5236 13962 5292 13972
rect 14522 13967 14532 14023
rect 14588 13967 14598 14023
rect 14746 13972 14756 14028
rect 14812 13972 14822 14028
rect 18788 13962 18844 13972
rect 18900 14028 18956 14038
rect 22820 14028 22876 14038
rect 19898 13972 19908 14028
rect 19964 13972 19974 14028
rect 22713 13977 22820 14023
rect 18900 13962 18956 13972
rect 22820 13962 22876 13972
rect 15988 13936 16044 13946
rect 4564 13916 4620 13926
rect 5796 13916 5852 13926
rect 7476 13916 7532 13926
rect 9716 13916 9772 13926
rect 2538 13860 2548 13916
rect 2604 13860 2614 13916
rect 3098 13860 3108 13916
rect 3164 13860 3174 13916
rect 3658 13860 3668 13916
rect 3724 13860 3734 13916
rect 3994 13860 4004 13916
rect 4060 13860 4070 13916
rect 4666 13860 4676 13916
rect 4732 13860 4742 13916
rect 6234 13860 6244 13916
rect 6300 13860 6310 13916
rect 7354 13860 7364 13916
rect 7420 13860 7430 13916
rect 7690 13860 7700 13916
rect 7756 13860 7766 13916
rect 9482 13860 9492 13916
rect 9548 13860 9558 13916
rect 4564 13850 4620 13860
rect 5796 13850 5852 13860
rect 7476 13850 7532 13860
rect 9716 13850 9772 13860
rect 10388 13916 10444 13926
rect 12068 13916 12124 13926
rect 10602 13860 10612 13916
rect 10668 13860 10678 13916
rect 13290 13860 13300 13916
rect 13356 13860 13366 13916
rect 15988 13870 16044 13880
rect 16436 13916 16492 13926
rect 22260 13916 22316 13926
rect 16538 13860 16548 13916
rect 16604 13860 16614 13916
rect 10388 13850 10444 13860
rect 12068 13850 12124 13860
rect 16436 13850 16492 13860
rect 22260 13850 22316 13860
rect 2996 13804 3052 13814
rect 12852 13804 12908 13814
rect 2996 13738 3052 13748
rect 6010 13692 6086 13738
rect 6010 13636 6020 13692
rect 6076 13636 6086 13692
rect 9370 13692 9446 13730
rect 9370 13636 9380 13692
rect 9436 13636 9446 13692
rect 10826 13692 10902 13792
rect 12852 13738 12908 13748
rect 17556 13804 17612 13814
rect 20794 13748 20804 13804
rect 20860 13748 20870 13804
rect 22138 13748 22148 13804
rect 22204 13748 22214 13804
rect 22922 13748 22932 13804
rect 22988 13748 22998 13804
rect 17556 13738 17612 13748
rect 10826 13636 10836 13692
rect 10892 13636 10902 13692
rect 16408 13468 16460 13524
rect 16516 13468 16616 13524
rect 16672 13468 16772 13524
rect 16828 13468 16928 13524
rect 16984 13468 17084 13524
rect 17140 13468 17192 13524
rect 1866 13300 1876 13356
rect 1932 13300 1942 13356
rect 2762 13300 2772 13356
rect 2828 13300 2838 13356
rect 3658 13300 3668 13356
rect 3724 13300 3734 13356
rect 4218 13300 4228 13356
rect 4284 13300 4294 13356
rect 1866 13262 1942 13300
rect 4218 13254 4294 13300
rect 11834 13300 11844 13356
rect 11900 13300 11910 13356
rect 11834 13254 11910 13300
rect 12954 13300 12964 13356
rect 13020 13300 13030 13356
rect 12954 13254 13030 13300
rect 19114 13300 19124 13356
rect 19180 13300 19190 13356
rect 19114 13262 19190 13300
rect 20570 13300 20580 13356
rect 20636 13300 20646 13356
rect 20570 13262 20646 13300
rect 1530 13239 1540 13244
rect 1402 13193 1540 13239
rect 1530 13188 1540 13193
rect 1596 13188 1606 13244
rect 9034 13188 9044 13244
rect 9100 13188 9110 13244
rect 18778 13239 18788 13244
rect 18650 13193 18788 13239
rect 18778 13188 18788 13193
rect 18844 13188 18854 13244
rect 196 13132 252 13142
rect 2212 13132 2268 13142
rect 3332 13132 3388 13142
rect 1082 13076 1092 13132
rect 1148 13076 1158 13132
rect 2314 13076 2324 13132
rect 2380 13076 2390 13132
rect 196 13066 252 13076
rect 2212 13066 2268 13076
rect 3332 13066 3388 13076
rect 3444 13132 3500 13142
rect 10500 13132 10556 13142
rect 4106 13076 4116 13132
rect 4172 13076 4182 13132
rect 4330 13076 4340 13132
rect 4396 13076 4406 13132
rect 4666 13076 4676 13132
rect 4732 13076 4742 13132
rect 8474 13076 8484 13132
rect 8540 13076 8550 13132
rect 3444 13066 3500 13076
rect 10500 13066 10556 13076
rect 11620 13132 11676 13142
rect 11620 13066 11676 13076
rect 12740 13132 12796 13142
rect 18116 13132 18172 13142
rect 14074 13076 14084 13132
rect 14140 13076 14150 13132
rect 12740 13066 12796 13076
rect 18116 13066 18172 13076
rect 19460 13132 19516 13142
rect 20132 13132 20188 13142
rect 19562 13076 19572 13132
rect 19628 13076 19638 13132
rect 19460 13066 19516 13076
rect 20132 13066 20188 13076
rect 20244 13132 20300 13142
rect 22148 13132 22204 13142
rect 21018 13076 21028 13132
rect 21084 13076 21094 13132
rect 21354 13076 21364 13132
rect 21420 13076 21430 13132
rect 20244 13066 20300 13076
rect 22148 13066 22204 13076
rect 22932 13132 22988 13142
rect 22932 13066 22988 13076
rect 12180 13020 12236 13030
rect 1754 12964 1764 13020
rect 1820 12964 1830 13020
rect 2426 12964 2436 13020
rect 2492 13015 2502 13020
rect 2492 12969 2599 13015
rect 2492 12964 2502 12969
rect 7130 12964 7140 13020
rect 7196 12964 7206 13020
rect 7354 12964 7364 13020
rect 7420 12964 7430 13020
rect 522 12908 598 12949
rect 4554 12908 4630 12949
rect 522 12852 532 12908
rect 588 12852 598 12908
rect 858 12852 868 12908
rect 924 12852 934 12908
rect 4554 12852 4564 12908
rect 4620 12852 4630 12908
rect 10042 12908 10118 13000
rect 11162 12964 11172 13020
rect 11228 12964 11238 13020
rect 15306 12964 15316 13020
rect 15372 12964 15382 13020
rect 15530 12964 15540 13020
rect 15596 12964 15606 13020
rect 17546 12964 17556 13020
rect 17612 12964 17622 13020
rect 18778 12964 18788 13020
rect 18844 13015 18854 13020
rect 18844 12969 19063 13015
rect 18844 12964 18854 12969
rect 20682 12964 20692 13020
rect 20748 12964 20758 13020
rect 21466 12969 21476 13025
rect 21532 12969 21542 13025
rect 12180 12954 12236 12964
rect 10042 12852 10052 12908
rect 10108 12852 10118 12908
rect 10714 12908 10790 12949
rect 22586 12908 22662 12949
rect 10714 12852 10724 12908
rect 10780 12852 10790 12908
rect 13402 12852 13412 12908
rect 13468 12903 13478 12908
rect 13468 12857 13687 12903
rect 13468 12852 13478 12857
rect 17994 12852 18004 12908
rect 18060 12852 18070 12908
rect 22586 12852 22596 12908
rect 22652 12852 22662 12908
rect 23258 12908 23334 12949
rect 23258 12852 23268 12908
rect 23324 12852 23334 12908
rect 10836 12796 10892 12806
rect 2986 12740 2996 12796
rect 3052 12740 3062 12796
rect 9818 12740 9828 12796
rect 9884 12740 9894 12796
rect 10836 12730 10892 12740
rect 11956 12796 12012 12806
rect 11956 12730 12012 12740
rect 5992 12572 6044 12628
rect 6100 12572 6200 12628
rect 6256 12572 6356 12628
rect 6412 12572 6512 12628
rect 6568 12572 6668 12628
rect 6724 12572 6776 12628
rect 5572 12460 5628 12470
rect 13748 12460 13804 12470
rect 4554 12404 4564 12460
rect 4620 12404 4630 12460
rect 13514 12404 13524 12460
rect 13580 12404 13590 12460
rect 5572 12394 5628 12404
rect 13748 12394 13804 12404
rect 14868 12460 14924 12470
rect 18218 12404 18228 12460
rect 18284 12404 18294 12460
rect 22922 12404 22932 12460
rect 22988 12455 22998 12460
rect 22988 12404 23110 12455
rect 14868 12394 14924 12404
rect 8820 12348 8876 12358
rect 6906 12343 6916 12348
rect 6249 12297 6916 12343
rect 6906 12292 6916 12297
rect 6972 12292 6982 12348
rect 8698 12343 8708 12348
rect 8586 12292 8708 12343
rect 8764 12292 8774 12348
rect 7588 12246 7644 12256
rect 4452 12236 4508 12246
rect 1082 12180 1092 12236
rect 1148 12180 1158 12236
rect 1306 12180 1316 12236
rect 1372 12180 1382 12236
rect 3546 12180 3556 12236
rect 3612 12231 3622 12236
rect 3612 12185 3719 12231
rect 3612 12180 3622 12185
rect 4452 12170 4508 12180
rect 7588 12170 7644 12190
rect 8026 12180 8036 12236
rect 8092 12180 8102 12236
rect 8362 12180 8372 12236
rect 8428 12180 8438 12236
rect 8586 12205 8662 12292
rect 8820 12282 8876 12292
rect 9604 12348 9660 12358
rect 23034 12356 23110 12404
rect 9604 12282 9660 12292
rect 12618 12292 12628 12348
rect 12684 12292 12694 12348
rect 12618 12251 12694 12292
rect 14746 12292 14756 12348
rect 14812 12292 14822 12348
rect 16874 12292 16884 12348
rect 16940 12343 16950 12348
rect 16940 12297 17398 12343
rect 16940 12292 16950 12297
rect 14746 12251 14822 12292
rect 17322 12251 17398 12297
rect 17994 12292 18004 12348
rect 18060 12292 18070 12348
rect 19114 12292 19124 12348
rect 19180 12292 19190 12348
rect 20122 12292 20132 12348
rect 20188 12292 20198 12348
rect 13412 12236 13468 12246
rect 15092 12236 15148 12246
rect 11274 12180 11284 12236
rect 11340 12180 11350 12236
rect 11498 12180 11508 12236
rect 11564 12180 11574 12236
rect 14074 12180 14084 12236
rect 14140 12180 14150 12236
rect 17994 12200 18070 12292
rect 20122 12251 20198 12292
rect 19786 12180 19796 12236
rect 19852 12231 19862 12236
rect 19852 12185 20071 12231
rect 19852 12180 19862 12185
rect 13412 12170 13468 12180
rect 15092 12170 15148 12180
rect 17556 12144 17612 12154
rect 3892 12124 3948 12134
rect 2426 12068 2436 12124
rect 2492 12068 2502 12124
rect 3210 12068 3220 12124
rect 3276 12068 3286 12124
rect 3892 12058 3948 12068
rect 5684 12124 5740 12134
rect 5684 12058 5740 12068
rect 5796 12124 5852 12134
rect 7466 12068 7476 12124
rect 7532 12068 7542 12124
rect 7802 12078 7812 12134
rect 7868 12078 7878 12134
rect 9044 12124 9100 12134
rect 8586 12068 8596 12124
rect 8652 12068 8662 12124
rect 5796 12058 5852 12068
rect 9044 12058 9100 12068
rect 9156 12124 9212 12134
rect 15876 12124 15932 12134
rect 10154 12068 10164 12124
rect 10220 12068 10230 12124
rect 12954 12068 12964 12124
rect 13020 12068 13030 12124
rect 14410 12068 14420 12124
rect 14476 12068 14486 12124
rect 15530 12068 15540 12124
rect 15596 12068 15606 12124
rect 19236 12124 19292 12134
rect 17556 12078 17612 12088
rect 18554 12068 18564 12124
rect 18620 12068 18630 12124
rect 9156 12058 9212 12068
rect 15876 12058 15932 12068
rect 19236 12058 19292 12068
rect 20468 12124 20524 12134
rect 20692 12124 20748 12134
rect 21924 12124 21980 12134
rect 20585 12073 20692 12119
rect 20468 12058 20524 12068
rect 21690 12068 21700 12124
rect 21756 12068 21766 12124
rect 20692 12058 20748 12068
rect 21924 12058 21980 12068
rect 22586 12063 22596 12119
rect 22652 12063 22662 12119
rect 5338 11956 5348 12012
rect 5404 12007 5414 12012
rect 5404 11961 5538 12007
rect 5404 11956 5414 11961
rect 7690 11956 7700 12012
rect 7756 11956 7766 12012
rect 7924 12007 7980 12017
rect 22820 12012 22876 12022
rect 19786 12007 19796 12012
rect 19658 11961 19796 12007
rect 19786 11956 19796 11961
rect 19852 11956 19862 12012
rect 21466 11956 21476 12012
rect 21532 11956 21558 12012
rect 7924 11941 7980 11951
rect 22820 11946 22876 11956
rect 6234 11900 6310 11938
rect 6234 11844 6244 11900
rect 6300 11844 6310 11900
rect 16408 11676 16460 11732
rect 16516 11676 16616 11732
rect 16672 11676 16772 11732
rect 16828 11676 16928 11732
rect 16984 11676 17084 11732
rect 17140 11676 17192 11732
rect 22148 11457 22204 11467
rect 5226 11396 5236 11452
rect 5292 11396 5302 11452
rect 21242 11396 21252 11452
rect 21308 11396 21318 11452
rect 22041 11401 22148 11447
rect 21242 11350 21318 11396
rect 22148 11391 22204 11401
rect 13748 11340 13804 11350
rect 20244 11340 20300 11350
rect 2986 11284 2996 11340
rect 3052 11284 3062 11340
rect 3994 11284 4004 11340
rect 4060 11335 4070 11340
rect 4330 11335 4340 11340
rect 4060 11289 4340 11335
rect 4060 11284 4070 11289
rect 4330 11284 4340 11289
rect 4396 11284 4406 11340
rect 4666 11284 4676 11340
rect 4732 11284 4742 11340
rect 7690 11284 7700 11340
rect 7756 11284 7766 11340
rect 12842 11284 12852 11340
rect 12908 11284 12918 11340
rect 17098 11284 17108 11340
rect 17164 11284 17174 11340
rect 13748 11274 13804 11284
rect 20244 11274 20300 11284
rect 21588 11340 21644 11350
rect 21588 11274 21644 11284
rect 22148 11335 22204 11345
rect 22204 11289 22311 11335
rect 22148 11269 22204 11279
rect 4564 11228 4620 11238
rect 13412 11228 13468 11238
rect 20020 11228 20076 11238
rect 22820 11228 22876 11238
rect 1642 11172 1652 11228
rect 1708 11172 1718 11228
rect 1866 11172 1876 11228
rect 1932 11172 1942 11228
rect 3770 11172 3780 11228
rect 3836 11172 3846 11228
rect 4793 11177 5002 11223
rect 6906 11172 6916 11228
rect 6972 11172 6982 11228
rect 8922 11172 8932 11228
rect 8988 11172 8998 11228
rect 9146 11172 9156 11228
rect 9212 11172 9222 11228
rect 11498 11172 11508 11228
rect 11564 11172 11574 11228
rect 11722 11172 11732 11228
rect 11788 11172 11798 11228
rect 14186 11172 14196 11228
rect 14252 11172 14262 11228
rect 16202 11172 16212 11228
rect 16268 11172 16278 11228
rect 18218 11172 18228 11228
rect 18284 11172 18294 11228
rect 18442 11172 18452 11228
rect 18508 11172 18518 11228
rect 20794 11172 20804 11228
rect 20860 11172 20870 11228
rect 22713 11177 22820 11223
rect 4564 11162 4620 11172
rect 13412 11162 13468 11172
rect 20020 11162 20076 11172
rect 22820 11162 22876 11172
rect 5226 11116 5302 11157
rect 5226 11060 5236 11116
rect 5292 11060 5302 11116
rect 13514 11116 13590 11157
rect 21018 11116 21094 11157
rect 13514 11060 13524 11116
rect 13580 11060 13590 11116
rect 19898 11060 19908 11116
rect 19964 11060 19974 11116
rect 21018 11060 21028 11116
rect 21084 11060 21094 11116
rect 23258 11060 23268 11116
rect 23324 11060 23370 11116
rect 14410 10948 14420 11004
rect 14476 10948 14486 11004
rect 5992 10780 6044 10836
rect 6100 10780 6200 10836
rect 6256 10780 6356 10836
rect 6412 10780 6512 10836
rect 6568 10780 6668 10836
rect 6724 10780 6776 10836
rect 12740 10668 12796 10678
rect 12740 10602 12796 10612
rect 13412 10668 13468 10678
rect 13412 10602 13468 10612
rect 15428 10556 15484 10566
rect 522 10500 532 10556
rect 588 10500 598 10556
rect 522 10459 598 10500
rect 11722 10500 11732 10556
rect 11788 10500 11798 10556
rect 11722 10459 11798 10500
rect 14522 10500 14532 10556
rect 14588 10500 14598 10556
rect 14522 10459 14598 10500
rect 15484 10505 15606 10551
rect 15428 10490 15484 10500
rect 15530 10459 15606 10505
rect 17434 10500 17444 10556
rect 17500 10551 17510 10556
rect 18666 10551 18676 10556
rect 17500 10505 17958 10551
rect 17500 10500 17510 10505
rect 17882 10459 17958 10505
rect 18554 10500 18676 10551
rect 18732 10500 18742 10556
rect 756 10444 812 10454
rect 11620 10444 11676 10454
rect 13636 10444 13692 10454
rect 18554 10450 18630 10500
rect 2742 10388 2752 10444
rect 2808 10388 2818 10444
rect 2986 10388 2996 10444
rect 3052 10388 3062 10444
rect 4106 10388 4116 10444
rect 4172 10388 4182 10444
rect 6010 10388 6020 10444
rect 6076 10388 6086 10444
rect 6234 10388 6244 10444
rect 6300 10388 6310 10444
rect 9706 10388 9716 10444
rect 9772 10388 9782 10444
rect 9930 10388 9940 10444
rect 9996 10388 10006 10444
rect 12394 10388 12404 10444
rect 12460 10388 12470 10444
rect 14298 10388 14308 10444
rect 14364 10388 14420 10444
rect 14858 10388 14868 10444
rect 14924 10388 14934 10444
rect 15866 10388 15876 10444
rect 15932 10388 15942 10444
rect 16202 10388 16212 10444
rect 16268 10388 16278 10444
rect 756 10378 812 10388
rect 11620 10378 11676 10388
rect 13636 10378 13692 10388
rect 196 10332 252 10342
rect 1204 10332 1260 10342
rect 970 10276 980 10332
rect 1036 10276 1046 10332
rect 196 10266 252 10276
rect 1204 10266 1260 10276
rect 1428 10332 1484 10342
rect 2324 10332 2380 10342
rect 1642 10276 1652 10332
rect 1708 10276 1718 10332
rect 3220 10332 3276 10342
rect 11956 10332 12012 10342
rect 2380 10281 2487 10327
rect 1428 10266 1484 10276
rect 2324 10266 2380 10276
rect 3322 10276 3332 10332
rect 3388 10276 3398 10332
rect 4778 10276 4788 10332
rect 4844 10276 4854 10332
rect 11050 10276 11060 10332
rect 11116 10276 11126 10332
rect 3220 10266 3276 10276
rect 3556 10220 3612 10230
rect 3408 10169 3556 10215
rect 3658 10220 3734 10270
rect 11956 10266 12012 10276
rect 14196 10332 14252 10342
rect 14196 10266 14252 10276
rect 15092 10332 15148 10342
rect 15092 10266 15148 10276
rect 15428 10332 15484 10342
rect 15428 10266 15484 10276
rect 15988 10332 16044 10342
rect 16202 10338 16278 10388
rect 18340 10439 18396 10449
rect 20020 10444 20076 10454
rect 19913 10393 20020 10439
rect 18340 10373 18396 10383
rect 20458 10388 20468 10444
rect 20524 10388 20534 10444
rect 22362 10388 22372 10444
rect 22428 10388 22438 10444
rect 22586 10388 22596 10444
rect 22652 10388 22662 10444
rect 20020 10378 20076 10388
rect 19348 10352 19404 10362
rect 15988 10266 16044 10276
rect 16324 10332 16380 10342
rect 16324 10266 16380 10276
rect 18228 10332 18284 10342
rect 19348 10286 19404 10296
rect 19460 10332 19516 10342
rect 18228 10266 18284 10276
rect 21130 10276 21140 10332
rect 21196 10276 21206 10332
rect 19460 10266 19516 10276
rect 3658 10164 3668 10220
rect 3724 10164 3734 10220
rect 19796 10220 19852 10230
rect 3556 10154 3612 10164
rect 1642 10108 1718 10154
rect 15204 10108 15270 10158
rect 19796 10154 19852 10164
rect 1642 10052 1652 10108
rect 1708 10052 1718 10108
rect 15194 10052 15204 10108
rect 15260 10052 15270 10108
rect 16408 9884 16460 9940
rect 16516 9884 16616 9940
rect 16672 9884 16772 9940
rect 16828 9884 16928 9940
rect 16984 9884 17084 9940
rect 17140 9884 17192 9940
rect 11844 9772 11900 9782
rect 634 9716 644 9772
rect 700 9716 710 9772
rect 970 9716 980 9772
rect 1036 9716 1046 9772
rect 634 9670 710 9716
rect 980 9666 1046 9716
rect 1306 9716 1316 9772
rect 1372 9716 1382 9772
rect 1306 9670 1382 9716
rect 11722 9716 11732 9772
rect 11788 9716 11798 9772
rect 11722 9670 11798 9716
rect 11900 9716 11910 9767
rect 11844 9670 11910 9716
rect 14746 9716 14756 9772
rect 14812 9716 14822 9772
rect 14746 9670 14822 9716
rect 14970 9716 14980 9772
rect 15036 9716 15046 9772
rect 14970 9660 15046 9716
rect 22474 9716 22484 9772
rect 22540 9716 22550 9772
rect 15988 9660 16044 9670
rect 10154 9604 10164 9660
rect 10220 9604 10230 9660
rect 22474 9622 22550 9716
rect 23706 9655 23716 9660
rect 23273 9609 23716 9655
rect 23706 9604 23716 9609
rect 23772 9604 23782 9660
rect 15988 9594 16044 9604
rect 74 9492 84 9548
rect 140 9492 150 9548
rect 746 9497 756 9553
rect 812 9497 822 9553
rect 1876 9548 1932 9558
rect 1194 9492 1204 9548
rect 1260 9492 1270 9548
rect 1540 9538 1596 9548
rect 1876 9482 1932 9492
rect 1988 9548 2044 9558
rect 2217 9497 2375 9543
rect 2650 9533 2660 9543
rect 1988 9482 2044 9492
rect 2553 9487 2660 9533
rect 2716 9487 2726 9543
rect 3882 9497 3892 9553
rect 3948 9497 3958 9553
rect 9268 9548 9324 9558
rect 10612 9548 10668 9558
rect 4106 9492 4116 9548
rect 4172 9492 4182 9548
rect 4666 9492 4676 9548
rect 4732 9492 4742 9548
rect 7914 9492 7924 9548
rect 7980 9492 7990 9548
rect 9818 9543 9828 9548
rect 9609 9497 9828 9543
rect 9818 9492 9828 9497
rect 9884 9492 9894 9548
rect 9268 9482 9324 9492
rect 10612 9482 10668 9492
rect 11508 9548 11564 9558
rect 13972 9548 14028 9558
rect 12170 9492 12180 9548
rect 12236 9492 12246 9548
rect 12954 9492 12964 9548
rect 13020 9543 13030 9548
rect 13020 9497 13127 9543
rect 13020 9492 13030 9497
rect 13738 9492 13748 9548
rect 13804 9492 13814 9548
rect 11508 9482 11564 9492
rect 13972 9482 14028 9492
rect 14084 9548 14140 9558
rect 14532 9548 14588 9558
rect 14186 9492 14196 9548
rect 14252 9492 14262 9548
rect 14634 9492 14644 9548
rect 14700 9492 14710 9548
rect 14858 9497 14868 9553
rect 14924 9497 14934 9553
rect 14980 9548 15036 9558
rect 15530 9502 15540 9558
rect 15596 9502 15606 9558
rect 15652 9548 15708 9558
rect 22260 9548 22316 9558
rect 14084 9482 14140 9492
rect 14532 9482 14588 9492
rect 14980 9482 15036 9492
rect 17098 9492 17108 9548
rect 17164 9543 17174 9548
rect 17164 9497 17271 9543
rect 17164 9492 17174 9497
rect 19674 9492 19684 9548
rect 19740 9492 19750 9548
rect 15652 9482 15708 9492
rect 22260 9482 22316 9492
rect 22932 9548 22988 9558
rect 22932 9482 22988 9492
rect 1540 9472 1596 9482
rect 3444 9436 3500 9446
rect 634 9370 644 9426
rect 700 9370 710 9426
rect 2650 9365 2660 9421
rect 2716 9375 2823 9421
rect 2716 9365 2726 9375
rect 3444 9370 3500 9380
rect 3668 9436 3724 9446
rect 9940 9436 9996 9446
rect 4228 9416 4284 9426
rect 3668 9370 3724 9380
rect 2314 9324 2390 9365
rect 3770 9355 3780 9411
rect 3836 9355 3846 9411
rect 6570 9380 6580 9436
rect 6636 9380 6646 9436
rect 6794 9380 6804 9436
rect 6860 9380 6870 9436
rect 8586 9380 8596 9436
rect 8652 9380 8662 9436
rect 9940 9370 9996 9380
rect 10948 9436 11004 9446
rect 10948 9370 11004 9380
rect 12628 9436 12684 9446
rect 17668 9436 17724 9446
rect 16090 9380 16100 9436
rect 16156 9380 16166 9436
rect 17892 9436 17948 9446
rect 17785 9385 17892 9431
rect 12628 9370 12684 9380
rect 4228 9350 4284 9360
rect 2314 9268 2324 9324
rect 2380 9268 2390 9324
rect 15306 9319 15382 9374
rect 17322 9324 17388 9374
rect 17668 9370 17724 9380
rect 18778 9380 18788 9436
rect 18844 9380 18854 9436
rect 20794 9380 20804 9436
rect 20860 9380 20870 9436
rect 21018 9380 21028 9436
rect 21084 9380 21094 9436
rect 17892 9370 17948 9380
rect 15530 9319 15540 9324
rect 15306 9273 15540 9319
rect 15530 9268 15540 9273
rect 15596 9268 15606 9324
rect 17322 9268 17332 9324
rect 17388 9268 17398 9324
rect 10724 9212 10780 9222
rect 12730 9156 12740 9212
rect 12796 9156 12806 9212
rect 10724 9146 10780 9156
rect 5992 8988 6044 9044
rect 6100 8988 6200 9044
rect 6256 8988 6356 9044
rect 6412 8988 6512 9044
rect 6568 8988 6668 9044
rect 6724 8988 6776 9044
rect 15428 8876 15484 8886
rect 1194 8820 1204 8876
rect 1260 8871 1270 8876
rect 1260 8825 1479 8871
rect 1260 8820 1270 8825
rect 1433 8759 1479 8825
rect 15428 8810 15484 8820
rect 1433 8713 2054 8759
rect 1978 8667 2054 8713
rect 2874 8708 2884 8764
rect 2940 8708 2950 8764
rect 5648 8708 5684 8764
rect 5740 8708 5750 8764
rect 7018 8708 7028 8764
rect 7084 8708 7094 8764
rect 8937 8713 9319 8759
rect 13626 8708 13636 8764
rect 13692 8759 13702 8764
rect 13692 8708 13814 8759
rect 2874 8658 2940 8708
rect 7018 8667 7094 8708
rect 13738 8667 13814 8708
rect 15306 8708 15316 8764
rect 15372 8708 15382 8764
rect 15306 8667 15382 8708
rect 16090 8708 16100 8764
rect 16156 8708 16166 8764
rect 9604 8652 9660 8662
rect 16090 8658 16166 8708
rect 16314 8708 16324 8764
rect 16380 8708 16390 8764
rect 16762 8708 16772 8764
rect 16828 8759 16838 8764
rect 17536 8759 17546 8764
rect 16828 8713 17286 8759
rect 16828 8708 16838 8713
rect 16314 8667 16390 8708
rect 17210 8667 17286 8713
rect 17434 8708 17546 8759
rect 17602 8708 17612 8764
rect 17882 8708 17892 8764
rect 17948 8708 17958 8764
rect 17434 8658 17510 8708
rect 17892 8667 17958 8708
rect 19226 8708 19236 8764
rect 19292 8708 19302 8764
rect 19562 8759 19572 8764
rect 298 8596 308 8652
rect 364 8596 374 8652
rect 970 8596 980 8652
rect 1036 8596 1046 8652
rect 2426 8596 2436 8652
rect 2492 8596 2502 8652
rect 2986 8596 2996 8652
rect 3052 8596 3062 8652
rect 3546 8596 3556 8652
rect 3612 8596 3622 8652
rect 11050 8596 11060 8652
rect 11116 8596 11126 8652
rect 11274 8596 11284 8652
rect 11340 8596 11350 8652
rect 13290 8596 13300 8652
rect 13356 8596 13366 8652
rect 17770 8596 17780 8652
rect 17836 8596 17846 8652
rect 19226 8621 19302 8708
rect 19460 8708 19572 8759
rect 19628 8708 19638 8764
rect 20122 8708 20132 8764
rect 20188 8708 20198 8764
rect 19460 8658 19526 8708
rect 20122 8667 20198 8708
rect 23482 8713 23492 8769
rect 23548 8713 23558 8769
rect 23482 8667 23558 8713
rect 20570 8647 20580 8652
rect 20473 8601 20580 8647
rect 20570 8596 20580 8601
rect 20636 8596 20646 8652
rect 308 8546 374 8596
rect 9604 8586 9660 8596
rect 2772 8540 2828 8550
rect 1082 8484 1092 8540
rect 1148 8484 1158 8540
rect 2650 8484 2660 8540
rect 2716 8484 2726 8540
rect 2772 8474 2828 8484
rect 3108 8540 3164 8550
rect 3892 8540 3948 8550
rect 3164 8489 3271 8535
rect 3322 8484 3332 8540
rect 3388 8484 3398 8540
rect 3770 8484 3780 8540
rect 3836 8484 3846 8540
rect 4106 8494 4116 8550
rect 4172 8494 4182 8550
rect 5460 8540 5516 8550
rect 5908 8540 5964 8550
rect 7252 8540 7308 8550
rect 8036 8540 8092 8550
rect 3108 8474 3164 8484
rect 3892 8474 3948 8484
rect 4340 8483 4396 8493
rect 84 8428 140 8438
rect 3434 8428 3510 8474
rect 3434 8372 3444 8428
rect 3500 8372 3510 8428
rect 5562 8484 5572 8540
rect 5628 8484 5638 8540
rect 5786 8484 5796 8540
rect 5852 8484 5862 8540
rect 6906 8484 6916 8540
rect 6972 8484 6982 8540
rect 7354 8484 7364 8540
rect 7420 8484 7430 8540
rect 7690 8484 7700 8540
rect 7756 8484 7766 8540
rect 4396 8432 4503 8478
rect 4340 8417 4396 8427
rect 5114 8428 5190 8478
rect 5460 8474 5516 8484
rect 5908 8474 5964 8484
rect 7252 8474 7308 8484
rect 8036 8474 8092 8484
rect 8148 8540 8204 8550
rect 9380 8540 9436 8550
rect 14644 8540 14700 8550
rect 8148 8474 8204 8484
rect 9268 8520 9324 8530
rect 12506 8484 12516 8540
rect 12572 8484 12582 8540
rect 14410 8484 14420 8540
rect 14476 8484 14486 8540
rect 14746 8484 14756 8540
rect 14812 8484 14822 8540
rect 15194 8484 15204 8540
rect 15260 8484 15270 8540
rect 15418 8484 15428 8540
rect 15484 8484 15494 8540
rect 15642 8489 15652 8545
rect 15708 8489 15718 8545
rect 15764 8540 15820 8550
rect 9380 8474 9436 8484
rect 14644 8474 14700 8484
rect 15764 8474 15820 8484
rect 18228 8540 18284 8550
rect 18676 8540 18732 8550
rect 18330 8484 18340 8540
rect 18396 8484 18406 8540
rect 18228 8474 18284 8484
rect 18676 8474 18732 8484
rect 19684 8540 19740 8550
rect 23044 8540 23100 8550
rect 20906 8484 20916 8540
rect 20972 8484 20982 8540
rect 19684 8474 19740 8484
rect 23044 8474 23100 8484
rect 9268 8454 9324 8464
rect 19124 8428 19180 8438
rect 5114 8372 5124 8428
rect 5180 8372 5190 8428
rect 7440 8372 7476 8428
rect 7532 8372 7542 8428
rect 14858 8372 14868 8428
rect 14924 8372 14934 8428
rect 16314 8372 16324 8428
rect 16380 8372 16390 8428
rect 17210 8372 17220 8428
rect 17276 8372 17286 8428
rect 84 8362 140 8372
rect 3556 8316 3622 8362
rect 3546 8260 3556 8316
rect 3612 8260 3622 8316
rect 4106 8316 4182 8372
rect 4106 8260 4116 8316
rect 4172 8260 4182 8316
rect 5450 8316 5526 8372
rect 5450 8260 5460 8316
rect 5516 8260 5526 8316
rect 7242 8316 7318 8372
rect 7242 8260 7252 8316
rect 7308 8260 7318 8316
rect 9706 8316 9782 8354
rect 9706 8260 9716 8316
rect 9772 8260 9782 8316
rect 18890 8316 18966 8410
rect 19180 8377 19287 8423
rect 22362 8372 22372 8428
rect 22428 8372 22438 8428
rect 19124 8362 19180 8372
rect 18890 8260 18900 8316
rect 18956 8260 18966 8316
rect 20682 8260 20692 8316
rect 20748 8260 20758 8316
rect 21466 8260 21476 8316
rect 21532 8260 21542 8316
rect 16408 8092 16460 8148
rect 16516 8092 16616 8148
rect 16672 8092 16772 8148
rect 16828 8092 16928 8148
rect 16984 8092 17084 8148
rect 17140 8092 17192 8148
rect 5562 7924 5572 7980
rect 5628 7924 5638 7980
rect 5562 7878 5638 7924
rect 9370 7924 9380 7980
rect 9436 7924 9446 7980
rect 9370 7878 9446 7924
rect 14410 7924 14420 7980
rect 14476 7924 14486 7980
rect 14410 7878 14486 7924
rect 14746 7924 14756 7980
rect 14812 7924 14822 7980
rect 15642 7924 15652 7980
rect 15708 7924 15718 7980
rect 14746 7874 14812 7924
rect 15642 7878 15718 7924
rect 16202 7924 16212 7980
rect 16268 7924 16278 7980
rect 16202 7868 16278 7924
rect 19684 7868 19740 7878
rect 17658 7812 17668 7868
rect 17724 7812 17734 7868
rect 19114 7812 19124 7868
rect 19180 7812 19190 7868
rect 17658 7802 17734 7812
rect 19684 7802 19740 7812
rect 21140 7868 21196 7878
rect 22138 7812 22148 7868
rect 22204 7863 22214 7868
rect 22204 7817 22342 7863
rect 22204 7812 22214 7817
rect 21140 7802 21196 7812
rect 4676 7756 4732 7766
rect 3210 7700 3220 7756
rect 3276 7700 3286 7756
rect 3994 7700 4004 7756
rect 4060 7700 4070 7756
rect 4442 7700 4452 7756
rect 4508 7700 4518 7756
rect 4676 7690 4732 7700
rect 4788 7756 4844 7766
rect 4788 7690 4844 7700
rect 5124 7756 5180 7766
rect 5796 7756 5852 7766
rect 5465 7705 5623 7751
rect 5124 7690 5180 7700
rect 5898 7700 5908 7756
rect 5964 7700 5974 7756
rect 6906 7705 6916 7761
rect 6972 7751 6982 7761
rect 9044 7756 9100 7766
rect 6972 7705 7191 7751
rect 7354 7700 7364 7756
rect 7420 7700 7430 7756
rect 7598 7700 7608 7756
rect 7664 7700 7674 7756
rect 5796 7690 5852 7700
rect 9044 7690 9100 7700
rect 9156 7756 9212 7766
rect 9156 7690 9212 7700
rect 9492 7756 9548 7766
rect 17658 7762 17724 7802
rect 18340 7756 18396 7766
rect 21476 7756 21532 7766
rect 13066 7700 13076 7756
rect 13132 7700 13142 7756
rect 14522 7700 14532 7756
rect 14588 7700 14598 7756
rect 14970 7700 14980 7756
rect 15036 7700 15046 7756
rect 15876 7736 15932 7746
rect 9492 7690 9548 7700
rect 15978 7700 15988 7756
rect 16044 7700 16054 7756
rect 16202 7700 16212 7756
rect 16268 7700 16278 7756
rect 16538 7700 16548 7756
rect 16604 7700 16614 7756
rect 17770 7700 17780 7756
rect 17836 7700 17846 7756
rect 18218 7700 18228 7756
rect 18284 7700 18294 7756
rect 19898 7700 19908 7756
rect 19964 7700 19974 7756
rect 21354 7700 21364 7756
rect 21420 7700 21430 7756
rect 15876 7670 15932 7680
rect 16100 7644 16156 7654
rect 1866 7588 1876 7644
rect 1932 7588 1942 7644
rect 2090 7588 2100 7644
rect 2156 7588 2166 7644
rect 10042 7639 10052 7644
rect 6906 7583 6916 7639
rect 6972 7583 6982 7639
rect 9945 7593 10052 7639
rect 10042 7588 10052 7593
rect 10108 7588 10118 7644
rect 11722 7588 11732 7644
rect 11788 7588 11798 7644
rect 11946 7588 11956 7644
rect 12012 7588 12022 7644
rect 15642 7588 15652 7644
rect 15708 7588 15718 7644
rect 16202 7639 16278 7700
rect 18340 7690 18396 7700
rect 21476 7690 21532 7700
rect 22708 7756 22764 7766
rect 22708 7690 22764 7700
rect 20916 7644 20972 7654
rect 16156 7593 16278 7639
rect 17434 7588 17444 7644
rect 17500 7588 17510 7644
rect 17994 7588 18004 7644
rect 18060 7588 18070 7644
rect 8250 7532 8326 7588
rect 16100 7578 16156 7588
rect 8250 7476 8260 7532
rect 8316 7476 8326 7532
rect 8698 7532 8774 7573
rect 8698 7476 8708 7532
rect 8764 7476 8774 7532
rect 13636 7532 13692 7542
rect 18666 7476 18676 7532
rect 18732 7527 18742 7532
rect 19114 7527 19190 7619
rect 19338 7588 19348 7644
rect 19404 7588 19414 7644
rect 20809 7593 20916 7639
rect 22138 7639 22148 7644
rect 21929 7593 22148 7639
rect 22138 7588 22148 7593
rect 22204 7588 22214 7644
rect 23370 7588 23380 7644
rect 23436 7588 23446 7644
rect 20916 7578 20972 7588
rect 21802 7532 21878 7573
rect 18732 7481 19190 7527
rect 18732 7476 18742 7481
rect 19562 7476 19572 7532
rect 19628 7527 19638 7532
rect 19628 7481 19735 7527
rect 19628 7476 19638 7481
rect 21802 7476 21812 7532
rect 21868 7476 21878 7532
rect 22922 7476 22932 7532
rect 22988 7476 22998 7532
rect 13636 7466 13692 7476
rect 17444 7420 17500 7430
rect 7354 7364 7364 7420
rect 7420 7364 7430 7420
rect 17444 7354 17500 7364
rect 18004 7420 18060 7430
rect 18004 7354 18060 7364
rect 5992 7196 6044 7252
rect 6100 7196 6200 7252
rect 6256 7196 6356 7252
rect 6412 7196 6512 7252
rect 6568 7196 6668 7252
rect 6724 7196 6776 7252
rect 14756 7084 14812 7094
rect 13178 7028 13188 7084
rect 13244 7028 13254 7084
rect 14756 7018 14812 7028
rect 12730 6916 12740 6972
rect 12796 6916 12806 6972
rect 12730 6875 12806 6916
rect 15642 6916 15652 6972
rect 15708 6916 15718 6972
rect 15642 6912 15718 6916
rect 15652 6875 15718 6912
rect 17770 6936 17780 6992
rect 17836 6936 17846 6992
rect 17770 6875 17836 6936
rect 19012 6880 19068 6890
rect 5796 6860 5852 6870
rect 1866 6804 1876 6860
rect 1932 6804 1942 6860
rect 2090 6804 2100 6860
rect 2156 6804 2166 6860
rect 3882 6804 3892 6860
rect 3948 6804 3958 6860
rect 6132 6860 6188 6870
rect 6025 6809 6132 6855
rect 5796 6794 5852 6804
rect 6132 6794 6188 6804
rect 7700 6860 7756 6870
rect 8586 6804 8596 6860
rect 8652 6804 8662 6860
rect 10602 6804 10612 6860
rect 10668 6804 10678 6860
rect 10826 6804 10836 6860
rect 10892 6804 10902 6860
rect 12506 6814 12516 6870
rect 12572 6814 12582 6870
rect 13300 6860 13356 6870
rect 7700 6794 7756 6804
rect 5236 6748 5292 6758
rect 5684 6748 5740 6758
rect 12506 6754 12572 6814
rect 13962 6804 13972 6860
rect 14028 6804 14084 6860
rect 14746 6804 14756 6860
rect 14812 6804 14822 6860
rect 16202 6819 16212 6875
rect 16268 6819 16278 6875
rect 18004 6870 18060 6880
rect 19012 6814 19068 6824
rect 19124 6865 19180 6875
rect 18004 6804 18060 6814
rect 13300 6794 13356 6804
rect 19124 6799 19180 6809
rect 22026 6804 22036 6860
rect 22092 6804 22102 6860
rect 13860 6748 13916 6758
rect 15092 6748 15148 6758
rect 15764 6748 15820 6758
rect 3210 6692 3220 6748
rect 3276 6692 3286 6748
rect 4666 6692 4676 6748
rect 4732 6692 4742 6748
rect 5114 6692 5124 6748
rect 5180 6692 5190 6748
rect 5450 6692 5460 6748
rect 5516 6743 5526 6748
rect 5516 6697 5623 6743
rect 5516 6692 5526 6697
rect 7802 6692 7812 6748
rect 7868 6692 7878 6748
rect 8250 6692 8260 6748
rect 8316 6692 8326 6748
rect 9482 6692 9492 6748
rect 9548 6692 9558 6748
rect 5236 6682 5292 6692
rect 5684 6682 5740 6692
rect 11946 6687 11956 6743
rect 12012 6687 12022 6743
rect 12618 6692 12628 6748
rect 12684 6692 12694 6748
rect 12954 6692 12964 6748
rect 13020 6692 13030 6748
rect 14970 6692 14980 6748
rect 15036 6692 15046 6748
rect 15530 6692 15540 6748
rect 15596 6692 15606 6748
rect 16314 6697 16324 6753
rect 16380 6697 16390 6753
rect 19908 6748 19964 6758
rect 17658 6692 17668 6748
rect 17724 6692 17734 6748
rect 17882 6692 17892 6748
rect 17948 6692 17958 6748
rect 19338 6692 19348 6748
rect 19404 6692 19414 6748
rect 19674 6692 19684 6748
rect 19740 6692 19750 6748
rect 13860 6682 13916 6692
rect 15092 6682 15148 6692
rect 15764 6682 15820 6692
rect 16650 6636 16726 6686
rect 15978 6580 15988 6636
rect 16044 6580 16054 6636
rect 16650 6580 16660 6636
rect 16716 6580 16726 6636
rect 18218 6636 18294 6686
rect 19908 6682 19964 6692
rect 20356 6748 20412 6758
rect 20356 6682 20412 6692
rect 20468 6748 20524 6758
rect 21028 6748 21084 6758
rect 20682 6692 20692 6748
rect 20748 6692 20758 6748
rect 21588 6748 21644 6758
rect 21257 6697 21527 6743
rect 20468 6682 20524 6692
rect 21028 6682 21084 6692
rect 21588 6682 21644 6692
rect 22820 6748 22876 6758
rect 23706 6743 23716 6748
rect 23273 6697 23716 6743
rect 23706 6692 23716 6697
rect 23772 6692 23782 6748
rect 22820 6682 22876 6692
rect 18218 6580 18228 6636
rect 18284 6580 18294 6636
rect 19226 6580 19236 6636
rect 19292 6580 19302 6636
rect 19424 6580 19460 6636
rect 19516 6580 19526 6636
rect 3770 6524 3846 6572
rect 3770 6468 3780 6524
rect 3836 6468 3846 6524
rect 4554 6524 4630 6570
rect 4554 6468 4564 6524
rect 4620 6468 4630 6524
rect 4890 6524 4956 6574
rect 8026 6524 8092 6574
rect 12506 6524 12582 6570
rect 4890 6468 4900 6524
rect 4956 6468 4966 6524
rect 8026 6468 8036 6524
rect 8092 6468 8102 6524
rect 12506 6468 12516 6524
rect 12572 6468 12582 6524
rect 16314 6514 16390 6575
rect 16314 6458 16324 6514
rect 16380 6458 16390 6514
rect 20010 6524 20086 6562
rect 20010 6468 20020 6524
rect 20076 6468 20086 6524
rect 21242 6524 21318 6570
rect 21242 6468 21252 6524
rect 21308 6468 21318 6524
rect 21914 6524 21990 6562
rect 21914 6468 21924 6524
rect 21980 6468 21990 6524
rect 16408 6300 16460 6356
rect 16516 6300 16616 6356
rect 16672 6300 16772 6356
rect 16828 6300 16928 6356
rect 16984 6300 17084 6356
rect 17140 6300 17192 6356
rect 4788 6188 4854 6199
rect 7476 6188 7532 6198
rect 4218 6132 4228 6188
rect 4284 6132 4294 6188
rect 4218 6086 4294 6132
rect 4788 6132 4798 6188
rect 5562 6132 5572 6188
rect 5628 6132 5638 6188
rect 4788 6082 4854 6132
rect 5572 6082 5638 6132
rect 6010 6132 6020 6188
rect 6076 6132 6086 6188
rect 6010 6086 6086 6132
rect 6906 6132 6916 6188
rect 6972 6132 6982 6188
rect 6906 6076 6982 6132
rect 7476 6122 7532 6132
rect 8036 6076 8092 6086
rect 3882 6020 3892 6076
rect 3948 6020 3958 6076
rect 5226 6020 5236 6076
rect 5292 6020 5302 6076
rect 7929 6025 8036 6071
rect 14176 6071 14186 6086
rect 14058 6030 14186 6071
rect 14242 6030 14252 6086
rect 14058 6025 14237 6030
rect 14522 6020 14532 6076
rect 14588 6020 14624 6076
rect 16650 6071 16660 6076
rect 16522 6025 16660 6071
rect 16650 6020 16660 6025
rect 16716 6020 16726 6076
rect 18554 6020 18564 6076
rect 18620 6020 18630 6076
rect 8036 6010 8092 6020
rect 20346 6015 20356 6071
rect 20412 6015 20422 6071
rect 4452 5964 4508 5974
rect 7588 5964 7644 5974
rect 12516 5969 12572 5979
rect 3098 5908 3108 5964
rect 3164 5908 3174 5964
rect 4452 5898 4508 5908
rect 4554 5903 4564 5959
rect 4620 5903 4630 5959
rect 5002 5908 5012 5964
rect 5068 5908 5078 5964
rect 5338 5908 5348 5964
rect 5404 5908 5414 5964
rect 5786 5908 5796 5964
rect 5852 5908 5862 5964
rect 6906 5908 6916 5964
rect 6972 5908 6982 5964
rect 7130 5908 7140 5964
rect 7196 5908 7252 5964
rect 7308 5908 7318 5964
rect 10490 5908 10500 5964
rect 10556 5908 10566 5964
rect 12394 5908 12404 5964
rect 12460 5908 12470 5964
rect 7588 5898 7644 5908
rect 12516 5903 12572 5913
rect 13636 5964 13692 5974
rect 16100 5964 16156 5974
rect 13636 5898 13692 5908
rect 14186 5903 14196 5959
rect 14252 5913 14359 5959
rect 14252 5903 14262 5913
rect 14634 5908 14644 5964
rect 14700 5908 14710 5964
rect 16100 5898 16156 5908
rect 17556 5964 17612 5974
rect 17556 5898 17612 5908
rect 19236 5964 19292 5974
rect 19338 5908 19348 5964
rect 19404 5908 19414 5964
rect 19236 5898 19292 5908
rect 1642 5796 1652 5852
rect 1708 5796 1718 5852
rect 1866 5796 1876 5852
rect 1932 5796 1942 5852
rect 7466 5740 7542 5827
rect 9146 5796 9156 5852
rect 9212 5796 9222 5852
rect 9370 5796 9380 5852
rect 9436 5796 9446 5852
rect 11274 5796 11284 5852
rect 11340 5796 11350 5852
rect 12730 5801 12740 5857
rect 12796 5801 12806 5857
rect 22260 5852 22316 5862
rect 12954 5796 12964 5852
rect 13020 5796 13030 5852
rect 15418 5796 15428 5852
rect 15484 5796 15494 5852
rect 18330 5796 18340 5852
rect 18396 5796 18406 5852
rect 18583 5827 18839 5847
rect 18554 5801 18839 5827
rect 21242 5796 21252 5852
rect 21308 5796 21318 5852
rect 22362 5796 22372 5852
rect 22428 5796 22438 5852
rect 22260 5786 22316 5796
rect 17994 5740 18070 5781
rect 7354 5684 7364 5740
rect 7420 5689 7542 5740
rect 12633 5735 12720 5740
rect 7420 5684 7430 5689
rect 12618 5679 12628 5735
rect 12684 5679 12720 5735
rect 13514 5684 13524 5740
rect 13580 5684 13590 5740
rect 15866 5684 15876 5740
rect 15932 5684 15942 5740
rect 17994 5684 18004 5740
rect 18060 5684 18070 5740
rect 18900 5715 18966 5781
rect 18890 5659 18900 5715
rect 18956 5659 18966 5715
rect 5992 5404 6044 5460
rect 6100 5404 6200 5460
rect 6256 5404 6356 5460
rect 6412 5404 6512 5460
rect 6568 5404 6668 5460
rect 6724 5404 6776 5460
rect 9706 5241 9716 5297
rect 9772 5241 9782 5297
rect 12628 5292 12684 5302
rect 11386 5236 11396 5292
rect 11452 5236 11462 5292
rect 12628 5226 12684 5236
rect 2314 5124 2324 5180
rect 2380 5124 2390 5180
rect 5114 5124 5124 5180
rect 5180 5124 5190 5180
rect 10154 5124 10164 5180
rect 10220 5175 10230 5180
rect 10220 5129 10566 5175
rect 10220 5124 10230 5129
rect 2324 5068 2390 5124
rect 4676 5078 4732 5088
rect 10490 5083 10566 5129
rect 12730 5124 12740 5180
rect 12796 5124 12806 5180
rect 12730 5083 12806 5124
rect 17770 5124 17780 5180
rect 17836 5124 17846 5180
rect 15652 5086 15708 5096
rect 17770 5087 17846 5124
rect 4004 5068 4060 5078
rect 2874 5012 2884 5068
rect 2940 5012 2950 5068
rect 3210 5012 3220 5068
rect 3276 5012 3286 5068
rect 4004 5002 4060 5012
rect 4116 5068 4172 5078
rect 4564 5068 4620 5078
rect 4172 5017 4391 5063
rect 4116 5002 4172 5012
rect 4900 5068 4956 5078
rect 4676 5012 4732 5022
rect 4793 5017 4900 5063
rect 11284 5068 11340 5078
rect 4564 5002 4620 5012
rect 4900 5002 4956 5012
rect 9604 5048 9660 5058
rect 11284 5002 11340 5012
rect 12404 5068 12460 5078
rect 12404 5002 12460 5012
rect 14644 5068 14700 5078
rect 15652 5020 15708 5030
rect 17210 5012 17220 5068
rect 17276 5012 17286 5068
rect 18666 5063 18676 5068
rect 18569 5017 18676 5063
rect 18666 5012 18676 5017
rect 18732 5012 18742 5068
rect 19002 5012 19012 5068
rect 19068 5012 19078 5068
rect 20346 5012 20356 5068
rect 20412 5012 20422 5068
rect 20570 5012 20580 5068
rect 20636 5012 20646 5068
rect 22474 5012 22484 5068
rect 22540 5012 22550 5068
rect 14644 5002 14700 5012
rect 9604 4982 9660 4992
rect 19002 4966 19078 5012
rect 1092 4956 1148 4966
rect 1764 4956 1820 4966
rect 74 4900 84 4956
rect 140 4900 150 4956
rect 410 4900 420 4956
rect 476 4900 486 4956
rect 1530 4900 1540 4956
rect 1596 4900 1606 4956
rect 1092 4890 1148 4900
rect 1764 4890 1820 4900
rect 1876 4956 1932 4966
rect 1876 4890 1932 4900
rect 2100 4956 2156 4966
rect 2436 4956 2492 4966
rect 2202 4900 2212 4956
rect 2268 4900 2278 4956
rect 2100 4890 2156 4900
rect 2436 4890 2492 4900
rect 2660 4956 2716 4966
rect 3444 4956 3500 4966
rect 2986 4900 2996 4956
rect 3052 4900 3062 4956
rect 3322 4900 3332 4956
rect 3388 4900 3398 4956
rect 2660 4890 2716 4900
rect 3444 4890 3500 4900
rect 3892 4956 3948 4966
rect 3892 4890 3948 4900
rect 5460 4956 5516 4966
rect 5684 4956 5740 4966
rect 5562 4900 5572 4956
rect 5628 4900 5638 4956
rect 5226 4844 5302 4894
rect 5460 4890 5516 4900
rect 5684 4890 5740 4900
rect 6132 4956 6188 4966
rect 8036 4956 8092 4966
rect 6346 4900 6356 4956
rect 6412 4900 6422 4956
rect 7242 4900 7252 4956
rect 7308 4900 7318 4956
rect 7593 4905 7751 4951
rect 6132 4890 6188 4900
rect 8036 4890 8092 4900
rect 8372 4956 8428 4966
rect 8596 4956 8652 4966
rect 12964 4956 13020 4966
rect 8474 4900 8484 4956
rect 8540 4900 8550 4956
rect 9146 4900 9156 4956
rect 9212 4900 9222 4956
rect 10826 4900 10836 4956
rect 10892 4900 10902 4956
rect 11946 4900 11956 4956
rect 12012 4900 12022 4956
rect 13402 4905 13412 4961
rect 13468 4905 13478 4961
rect 13636 4956 13692 4966
rect 13972 4956 14028 4966
rect 8372 4890 8428 4900
rect 8596 4890 8652 4900
rect 12964 4890 13020 4900
rect 13850 4900 13860 4956
rect 13916 4900 13926 4956
rect 14868 4956 14924 4966
rect 15764 4956 15820 4966
rect 14089 4905 14471 4951
rect 13636 4890 13692 4900
rect 13972 4890 14028 4900
rect 15301 4900 15311 4956
rect 15367 4900 15377 4956
rect 14868 4890 14924 4900
rect 15530 4890 15540 4946
rect 15596 4890 15606 4946
rect 15764 4890 15820 4900
rect 17556 4956 17612 4966
rect 18116 4956 18172 4966
rect 22932 4956 22988 4966
rect 17785 4905 18055 4951
rect 17556 4890 17612 4900
rect 21690 4900 21700 4956
rect 21756 4900 21766 4956
rect 23706 4951 23716 4956
rect 23385 4905 23716 4951
rect 23706 4900 23716 4905
rect 23772 4900 23782 4956
rect 18116 4890 18172 4900
rect 22932 4890 22988 4900
rect 6244 4844 6300 4854
rect 5226 4788 5236 4844
rect 5292 4788 5302 4844
rect 5898 4788 5908 4844
rect 5964 4788 5974 4844
rect 7466 4788 7476 4844
rect 7532 4788 7568 4844
rect 14298 4839 14308 4844
rect 14062 4793 14308 4839
rect 14298 4788 14308 4793
rect 14364 4788 14374 4844
rect 74 4732 150 4788
rect 2650 4732 2726 4782
rect 6244 4778 6300 4788
rect 74 4676 84 4732
rect 140 4676 150 4732
rect 2538 4676 2548 4732
rect 2604 4681 2726 4732
rect 3658 4732 3734 4778
rect 2604 4676 2614 4681
rect 3658 4676 3668 4732
rect 3724 4676 3734 4732
rect 8810 4732 8886 4778
rect 8810 4676 8820 4732
rect 8876 4676 8886 4732
rect 11610 4732 11686 4778
rect 11610 4676 11620 4732
rect 11676 4676 11686 4732
rect 18442 4732 18518 4770
rect 18442 4676 18452 4732
rect 18508 4676 18518 4732
rect 18778 4732 18854 4778
rect 18778 4676 18788 4732
rect 18844 4676 18854 4732
rect 16408 4508 16460 4564
rect 16516 4508 16616 4564
rect 16672 4508 16772 4564
rect 16828 4508 16928 4564
rect 16984 4508 17084 4564
rect 17140 4508 17192 4564
rect 858 4340 868 4396
rect 924 4340 934 4396
rect 308 4284 364 4294
rect 858 4293 934 4340
rect 2874 4340 2884 4396
rect 2940 4340 2950 4396
rect 4106 4345 4116 4401
rect 4172 4345 4182 4401
rect 2874 4290 2940 4340
rect 4106 4294 4182 4345
rect 4442 4340 4452 4396
rect 4508 4340 4518 4396
rect 4442 4294 4518 4340
rect 13402 4340 13412 4396
rect 13468 4340 13478 4396
rect 13402 4292 13478 4340
rect 15418 4340 15428 4396
rect 15484 4340 15494 4396
rect 15418 4294 15494 4340
rect 2426 4228 2436 4284
rect 2492 4228 2502 4284
rect 4778 4228 4788 4284
rect 4844 4228 4880 4284
rect 17870 4228 17892 4284
rect 17948 4228 17958 4284
rect 23482 4279 23492 4284
rect 23385 4233 23492 4279
rect 23482 4228 23492 4233
rect 23548 4228 23558 4284
rect 308 4218 364 4228
rect 84 4172 140 4182
rect 84 4106 140 4116
rect 420 4172 476 4182
rect 420 4106 476 4116
rect 980 4172 1036 4182
rect 1540 4172 1596 4182
rect 1876 4172 1932 4182
rect 1306 4116 1316 4172
rect 1372 4116 1382 4172
rect 1642 4116 1652 4172
rect 1708 4116 1718 4172
rect 980 4106 1036 4116
rect 1540 4106 1596 4116
rect 1876 4106 1932 4116
rect 1988 4172 2044 4182
rect 14308 4172 14364 4182
rect 17444 4172 17500 4182
rect 23044 4172 23100 4182
rect 2314 4116 2324 4172
rect 2380 4116 2390 4172
rect 2650 4116 2660 4172
rect 2716 4116 2726 4172
rect 3098 4116 3108 4172
rect 3164 4116 3174 4172
rect 3770 4116 3780 4172
rect 3836 4116 3846 4172
rect 4106 4116 4116 4172
rect 4172 4116 4182 4172
rect 4330 4116 4340 4172
rect 4396 4116 4406 4172
rect 4554 4116 4564 4172
rect 4620 4116 4630 4172
rect 4890 4116 4900 4172
rect 4956 4116 4966 4172
rect 8698 4116 8708 4172
rect 8764 4116 8774 4172
rect 12842 4116 12852 4172
rect 12908 4116 12918 4172
rect 14858 4116 14868 4172
rect 14924 4116 14934 4172
rect 16986 4116 16996 4172
rect 17052 4116 17062 4172
rect 18330 4116 18340 4172
rect 18396 4116 18406 4172
rect 18778 4116 18788 4172
rect 18844 4116 18854 4172
rect 22138 4116 22148 4172
rect 22204 4167 22214 4172
rect 22204 4121 22311 4167
rect 22204 4116 22214 4121
rect 1988 4106 2044 4116
rect 14308 4106 14364 4116
rect 23044 4106 23100 4116
rect 2212 4060 2268 4070
rect 7354 4004 7364 4060
rect 7420 4004 7430 4060
rect 7578 4004 7588 4060
rect 7644 4004 7654 4060
rect 9594 4004 9604 4060
rect 9660 4004 9670 4060
rect 11498 4004 11508 4060
rect 11564 4004 11574 4060
rect 11722 4004 11732 4060
rect 11788 4004 11798 4060
rect 14074 4055 14150 4094
rect 13852 4009 14150 4055
rect 14420 4060 14476 4070
rect 20020 4060 20076 4070
rect 21588 4060 21644 4070
rect 15158 4004 15204 4060
rect 15260 4004 15270 4060
rect 17882 4004 17892 4060
rect 17948 4055 17958 4060
rect 17948 4009 18167 4055
rect 17948 4004 17958 4009
rect 19898 4004 19908 4060
rect 19964 4004 19974 4060
rect 21018 4004 21028 4060
rect 21084 4004 21094 4060
rect 22820 4060 22876 4070
rect 22713 4009 22820 4055
rect 2212 3994 2268 4004
rect 14420 3994 14476 4004
rect 14746 3948 14822 3989
rect 18554 3948 18620 3998
rect 20020 3994 20076 4004
rect 21588 3994 21644 4004
rect 22820 3994 22876 4004
rect 14746 3892 14756 3948
rect 14812 3892 14822 3948
rect 17210 3892 17220 3948
rect 17276 3892 17286 3948
rect 18554 3892 18564 3948
rect 18620 3892 18630 3948
rect 17780 3836 17836 3846
rect 17780 3770 17836 3780
rect 5992 3612 6044 3668
rect 6100 3612 6200 3668
rect 6256 3612 6356 3668
rect 6412 3612 6512 3668
rect 6568 3612 6668 3668
rect 6724 3612 6776 3668
rect 13636 3500 13692 3510
rect 4554 3444 4564 3500
rect 4620 3444 4712 3500
rect 5002 3444 5012 3500
rect 5068 3444 5078 3500
rect 1418 3332 1428 3388
rect 1484 3332 1494 3388
rect 4442 3337 4452 3393
rect 4508 3383 4518 3393
rect 5786 3388 5862 3444
rect 13636 3434 13692 3444
rect 4508 3337 4630 3383
rect 3444 3276 3500 3286
rect 4554 3276 4630 3337
rect 5786 3332 5796 3388
rect 5852 3332 5862 3388
rect 13290 3332 13300 3388
rect 13356 3332 13366 3388
rect 12516 3276 12572 3286
rect 858 3220 868 3276
rect 924 3220 934 3276
rect 1530 3220 1540 3276
rect 1596 3220 1606 3276
rect 2202 3220 2212 3276
rect 2268 3220 2278 3276
rect 8250 3220 8260 3276
rect 8316 3220 8326 3276
rect 858 3216 934 3220
rect 868 3170 934 3216
rect 3444 3210 3500 3220
rect 10042 3215 10052 3271
rect 10108 3215 10118 3271
rect 10266 3220 10276 3276
rect 10332 3220 10342 3276
rect 12572 3225 12679 3271
rect 13290 3240 13366 3332
rect 13850 3332 13860 3388
rect 13916 3332 13926 3388
rect 13850 3291 13926 3332
rect 15306 3332 15316 3388
rect 15372 3332 15382 3388
rect 15306 3282 15382 3332
rect 15978 3332 15988 3388
rect 16044 3332 16054 3388
rect 15978 3291 16054 3332
rect 17210 3332 17220 3388
rect 17276 3332 17286 3388
rect 20234 3332 20244 3388
rect 20300 3332 20310 3388
rect 17210 3322 17286 3332
rect 17220 3282 17286 3322
rect 20244 3282 20310 3332
rect 23034 3332 23044 3388
rect 23100 3332 23110 3388
rect 23034 3291 23110 3332
rect 21476 3276 21532 3286
rect 15082 3220 15092 3276
rect 15148 3220 15158 3276
rect 17434 3220 17444 3276
rect 17500 3220 17556 3276
rect 17770 3220 17780 3276
rect 17836 3220 17882 3276
rect 18518 3220 18564 3276
rect 18620 3220 18630 3276
rect 19002 3220 19012 3276
rect 19068 3220 19114 3276
rect 20794 3220 20804 3276
rect 20860 3220 20906 3276
rect 21466 3220 21476 3271
rect 21588 3276 21644 3286
rect 21532 3220 21542 3271
rect 12516 3210 12572 3220
rect 21466 3174 21542 3220
rect 21924 3276 21980 3286
rect 21588 3210 21644 3220
rect 21802 3225 21924 3271
rect 21802 3174 21878 3225
rect 21924 3210 21980 3220
rect 23380 3276 23436 3286
rect 23380 3210 23436 3220
rect 2436 3164 2492 3174
rect 2436 3098 2492 3108
rect 2548 3164 2604 3174
rect 2548 3098 2604 3108
rect 2772 3164 2828 3174
rect 2772 3098 2828 3108
rect 3780 3164 3836 3174
rect 4116 3164 4172 3174
rect 5460 3164 5516 3174
rect 7924 3164 7980 3174
rect 8708 3164 8764 3174
rect 3882 3108 3892 3164
rect 3948 3108 3958 3164
rect 4218 3108 4228 3164
rect 4284 3108 4294 3164
rect 4554 3159 4564 3164
rect 4457 3113 4564 3159
rect 4554 3108 4564 3113
rect 4620 3108 4630 3164
rect 5226 3108 5236 3164
rect 5292 3108 5302 3164
rect 7354 3108 7364 3164
rect 7420 3108 7430 3164
rect 7690 3108 7700 3164
rect 7756 3108 7766 3164
rect 8026 3108 8036 3164
rect 8092 3108 8102 3164
rect 3780 3098 3836 3108
rect 4116 3098 4172 3108
rect 5460 3098 5516 3108
rect 7924 3098 7980 3108
rect 8708 3098 8764 3108
rect 8820 3164 8876 3174
rect 18228 3164 18284 3174
rect 22484 3164 22540 3174
rect 11498 3108 11508 3164
rect 11564 3108 11574 3164
rect 12954 3108 12964 3164
rect 13020 3108 13030 3164
rect 14074 3108 14084 3164
rect 14140 3108 14150 3164
rect 8820 3098 8876 3108
rect 14746 3103 14756 3159
rect 14812 3103 14822 3159
rect 15306 3108 15316 3164
rect 15372 3108 15382 3164
rect 15642 3108 15652 3164
rect 15708 3159 15718 3164
rect 15708 3113 15815 3159
rect 15708 3108 15718 3113
rect 16090 3108 16100 3164
rect 16156 3108 16166 3164
rect 16986 3108 16996 3164
rect 17052 3108 17062 3164
rect 18106 3108 18116 3164
rect 18172 3108 18182 3164
rect 19338 3108 19348 3164
rect 19404 3108 19414 3164
rect 20010 3108 20020 3164
rect 20076 3108 20086 3164
rect 21145 3113 21303 3159
rect 644 3052 700 3062
rect 14634 3052 14700 3102
rect 18228 3098 18284 3108
rect 22484 3098 22540 3108
rect 22596 3164 22652 3174
rect 22596 3098 22652 3108
rect 8586 2996 8596 3052
rect 8652 2996 8662 3052
rect 12282 2996 12292 3052
rect 12348 2996 12358 3052
rect 14634 2996 14644 3052
rect 14700 2996 14710 3052
rect 644 2986 700 2996
rect 1866 2940 1942 2987
rect 7690 2940 7766 2986
rect 1866 2884 1876 2940
rect 1932 2884 1942 2940
rect 4778 2884 4788 2940
rect 4844 2884 4854 2940
rect 7690 2884 7700 2940
rect 7756 2884 7766 2940
rect 8250 2940 8326 2986
rect 8250 2884 8260 2940
rect 8316 2884 8326 2940
rect 18778 2940 18854 2978
rect 18778 2884 18788 2940
rect 18844 2884 18854 2940
rect 20570 2940 20646 2978
rect 20570 2884 20580 2940
rect 20636 2884 20646 2940
rect 22138 2940 22214 3034
rect 22138 2884 22148 2940
rect 22204 2884 22214 2940
rect 16408 2716 16460 2772
rect 16516 2716 16616 2772
rect 16672 2716 16772 2772
rect 16828 2716 16928 2772
rect 16984 2716 17084 2772
rect 17140 2716 17192 2772
rect 4218 2548 4228 2604
rect 4284 2548 4294 2604
rect 4218 2502 4294 2548
rect 7466 2548 7476 2604
rect 7532 2548 7542 2604
rect 3882 2436 3892 2492
rect 3948 2436 3958 2492
rect 5114 2436 5124 2492
rect 5180 2436 5206 2492
rect 7466 2464 7542 2548
rect 9258 2548 9268 2604
rect 9324 2548 9334 2604
rect 9930 2548 9940 2604
rect 9996 2548 10006 2604
rect 9258 2492 9334 2548
rect 9940 2498 10006 2548
rect 15642 2548 15652 2604
rect 15708 2548 15718 2604
rect 15642 2502 15718 2548
rect 18218 2548 18228 2604
rect 18284 2548 18294 2604
rect 18218 2502 18294 2548
rect 18666 2548 18676 2604
rect 18732 2548 18742 2604
rect 18666 2502 18742 2548
rect 18004 2492 18060 2502
rect 10378 2436 10388 2492
rect 10444 2436 10454 2492
rect 17897 2441 18004 2487
rect 18004 2426 18060 2436
rect 5572 2380 5628 2390
rect 8708 2380 8764 2390
rect 9156 2380 9212 2390
rect 9604 2380 9660 2390
rect 14532 2380 14588 2390
rect 3098 2324 3108 2380
rect 3164 2324 3174 2380
rect 4442 2324 4452 2380
rect 4508 2324 4518 2380
rect 4905 2329 5063 2375
rect 1642 2212 1652 2268
rect 1708 2212 1718 2268
rect 1866 2212 1876 2268
rect 1932 2212 1942 2268
rect 5017 2263 5063 2329
rect 5572 2314 5628 2324
rect 7690 2319 7700 2375
rect 7756 2319 7766 2375
rect 8586 2324 8596 2380
rect 8652 2324 8662 2380
rect 8922 2324 8932 2380
rect 8988 2324 8998 2380
rect 9258 2324 9268 2380
rect 9324 2324 9334 2380
rect 9706 2324 9716 2380
rect 9772 2324 9782 2380
rect 10154 2324 10164 2380
rect 10220 2324 10230 2380
rect 10490 2324 10500 2380
rect 10556 2324 10566 2380
rect 10826 2324 10836 2380
rect 10892 2324 10902 2380
rect 11050 2324 11060 2380
rect 11116 2324 11126 2380
rect 11722 2324 11732 2380
rect 11788 2324 11798 2380
rect 12282 2324 12292 2380
rect 12348 2324 12358 2380
rect 13178 2324 13188 2380
rect 13244 2324 13290 2380
rect 13514 2324 13524 2380
rect 13580 2324 13590 2380
rect 14186 2324 14196 2380
rect 14252 2324 14262 2380
rect 8708 2314 8764 2324
rect 9156 2314 9212 2324
rect 9604 2314 9660 2324
rect 14532 2314 14588 2324
rect 14644 2380 14700 2390
rect 14644 2314 14700 2324
rect 14858 2380 14914 2390
rect 14858 2314 14914 2324
rect 14980 2380 15036 2390
rect 14980 2314 15036 2324
rect 15316 2380 15372 2390
rect 15316 2314 15372 2324
rect 15876 2380 15932 2390
rect 16548 2380 16604 2390
rect 18116 2380 18172 2390
rect 15978 2324 15988 2380
rect 16044 2324 16054 2380
rect 16202 2324 16212 2380
rect 16268 2324 16278 2380
rect 16426 2324 16436 2380
rect 16492 2324 16502 2380
rect 16762 2324 16772 2380
rect 16828 2324 16838 2380
rect 15876 2314 15932 2324
rect 16548 2314 16604 2324
rect 18116 2314 18172 2324
rect 18340 2380 18396 2390
rect 18340 2314 18396 2324
rect 18452 2380 18508 2390
rect 18452 2314 18508 2324
rect 18788 2380 18844 2390
rect 21018 2324 21028 2380
rect 21084 2324 21094 2380
rect 21130 2324 21140 2380
rect 21196 2324 21206 2380
rect 18788 2314 18844 2324
rect 5114 2263 5124 2268
rect 5017 2217 5124 2263
rect 5114 2212 5124 2217
rect 5180 2212 5190 2268
rect 6234 2212 6244 2268
rect 6300 2212 6310 2268
rect 3658 2156 3734 2197
rect 3658 2100 3668 2156
rect 3724 2100 3734 2156
rect 4666 2166 4732 2206
rect 8026 2202 8036 2258
rect 8092 2202 8102 2258
rect 11162 2212 11172 2268
rect 11228 2212 11238 2268
rect 14410 2212 14420 2268
rect 14476 2212 14486 2268
rect 17658 2212 17668 2268
rect 17724 2212 17734 2268
rect 4666 2156 4742 2166
rect 4666 2100 4676 2156
rect 4732 2100 4742 2156
rect 5338 2100 5348 2156
rect 5404 2100 5414 2156
rect 8250 2151 8326 2197
rect 8250 2095 8260 2151
rect 8316 2095 8326 2151
rect 10602 2156 10678 2197
rect 10602 2100 10612 2156
rect 10668 2100 10678 2156
rect 13514 2146 13590 2197
rect 15204 2156 15270 2206
rect 19114 2156 19190 2243
rect 20346 2212 20356 2268
rect 20412 2212 20422 2268
rect 22250 2212 22260 2268
rect 22316 2212 22326 2268
rect 22474 2212 22484 2268
rect 22540 2212 22550 2268
rect 13514 2090 13524 2146
rect 13580 2090 13590 2146
rect 15194 2100 15204 2156
rect 15260 2100 15270 2156
rect 15642 2100 15652 2156
rect 15708 2151 15718 2156
rect 15708 2105 15927 2151
rect 15708 2100 15718 2105
rect 19114 2100 19124 2156
rect 19180 2100 19190 2156
rect 16772 2044 16828 2054
rect 16772 1978 16828 1988
rect 5992 1820 6044 1876
rect 6100 1820 6200 1876
rect 6256 1820 6356 1876
rect 6412 1820 6512 1876
rect 6568 1820 6668 1876
rect 6724 1820 6776 1876
rect 17556 1708 17612 1718
rect 17556 1642 17612 1652
rect 2314 1540 2324 1596
rect 2380 1540 2390 1596
rect 3546 1540 3556 1596
rect 3612 1540 3622 1596
rect 4218 1540 4228 1596
rect 4284 1540 4294 1596
rect 4218 1499 4294 1540
rect 5114 1540 5124 1596
rect 5180 1540 5190 1596
rect 5562 1540 5572 1596
rect 5628 1540 5638 1596
rect 7690 1540 7700 1596
rect 7756 1540 7766 1596
rect 9930 1540 9940 1596
rect 9996 1540 10006 1596
rect 13290 1540 13300 1596
rect 13356 1540 13366 1596
rect 5114 1499 5190 1540
rect 13290 1499 13366 1540
rect 13962 1540 13972 1596
rect 14028 1540 14038 1596
rect 13962 1499 14038 1540
rect 14522 1540 14532 1596
rect 14588 1540 14598 1596
rect 1204 1484 1260 1494
rect 14522 1484 14598 1540
rect 14746 1540 14756 1596
rect 14812 1540 14822 1596
rect 17098 1591 17108 1596
rect 14746 1530 14822 1540
rect 16650 1545 17108 1591
rect 14746 1490 14812 1530
rect 16650 1499 16726 1545
rect 17098 1540 17108 1545
rect 17164 1540 17174 1596
rect 15316 1484 15372 1494
rect 298 1428 308 1484
rect 364 1428 374 1484
rect 858 1428 868 1484
rect 924 1428 934 1484
rect 1204 1418 1260 1428
rect 1754 1428 1764 1484
rect 1820 1428 1830 1484
rect 2426 1428 2436 1484
rect 2492 1428 2502 1484
rect 2986 1428 2996 1484
rect 3052 1428 3062 1484
rect 3658 1428 3668 1484
rect 3724 1428 3734 1484
rect 7578 1428 7588 1484
rect 7644 1428 7654 1484
rect 1754 1424 1830 1428
rect 2986 1424 3062 1428
rect 1764 1378 1830 1424
rect 2772 1372 2828 1382
rect 2996 1378 3062 1424
rect 15316 1418 15372 1428
rect 16212 1479 16268 1489
rect 16212 1413 16268 1423
rect 16324 1479 16380 1489
rect 18564 1484 18620 1494
rect 17882 1428 17892 1484
rect 17948 1428 17958 1484
rect 20234 1428 20244 1484
rect 20300 1428 20310 1484
rect 20458 1428 20468 1484
rect 20524 1428 20534 1484
rect 22250 1428 22260 1484
rect 22316 1428 22326 1484
rect 16324 1413 16380 1423
rect 18564 1418 18620 1428
rect 12068 1372 12124 1382
rect 15092 1372 15148 1382
rect 186 1316 196 1372
rect 252 1316 262 1372
rect 1433 1321 1591 1367
rect 3994 1316 4004 1372
rect 4060 1316 4070 1372
rect 4330 1316 4340 1372
rect 4396 1316 4406 1372
rect 5002 1316 5012 1372
rect 5068 1316 5078 1372
rect 5353 1321 5572 1367
rect 5674 1316 5684 1372
rect 5740 1316 5750 1372
rect 6010 1316 6020 1372
rect 6076 1316 6086 1372
rect 6346 1316 6356 1372
rect 6412 1316 6422 1372
rect 8138 1316 8148 1372
rect 8204 1316 8214 1372
rect 9818 1316 9828 1372
rect 9884 1316 9894 1372
rect 10378 1316 10388 1372
rect 10444 1316 10454 1372
rect 11386 1367 11396 1372
rect 11042 1321 11396 1367
rect 11386 1316 11396 1321
rect 11452 1316 11462 1372
rect 12282 1316 12292 1372
rect 12348 1316 12358 1372
rect 12730 1316 12740 1372
rect 12796 1316 12806 1372
rect 13030 1316 13076 1372
rect 13132 1316 13142 1372
rect 2772 1306 2828 1316
rect 12068 1306 12124 1316
rect 13402 1311 13412 1367
rect 13468 1311 13478 1367
rect 13702 1316 13748 1372
rect 13804 1316 13814 1372
rect 14522 1316 14532 1372
rect 14588 1316 14598 1372
rect 14970 1316 14980 1372
rect 15036 1316 15046 1372
rect 15092 1306 15148 1316
rect 15978 1311 15988 1367
rect 16044 1311 16054 1367
rect 18218 1316 18228 1372
rect 18284 1316 18294 1372
rect 21578 1316 21588 1372
rect 21644 1316 21654 1372
rect 23706 1367 23716 1372
rect 22438 1321 22871 1367
rect 23273 1321 23716 1367
rect 23706 1316 23716 1321
rect 23772 1316 23782 1372
rect 8698 1204 8708 1260
rect 8764 1204 8774 1260
rect 12618 1255 12628 1260
rect 12490 1209 12628 1255
rect 12618 1204 12628 1209
rect 12684 1204 12694 1260
rect 16408 924 16460 980
rect 16516 924 16616 980
rect 16672 924 16772 980
rect 16828 924 16928 980
rect 16984 924 17084 980
rect 17140 924 17192 980
rect 4442 756 4452 812
rect 4508 756 4518 812
rect 12170 756 12180 812
rect 12236 756 12246 812
rect 15754 756 15764 812
rect 15820 756 15830 812
rect 4442 664 4518 756
rect 15754 718 15830 756
rect 9258 644 9268 700
rect 9324 644 9334 700
rect 20682 644 20692 700
rect 20748 644 20758 700
rect 4900 588 4956 598
rect 10500 588 10556 598
rect 3098 532 3108 588
rect 3164 532 3174 588
rect 4666 532 4676 588
rect 4732 532 4742 588
rect 8698 532 8708 588
rect 8764 532 8774 588
rect 4900 522 4956 532
rect 10500 522 10556 532
rect 11508 588 11564 598
rect 13412 588 13468 598
rect 15092 588 15148 598
rect 12842 532 12852 588
rect 12908 532 12918 588
rect 13514 532 13524 588
rect 13580 532 13590 588
rect 14074 532 14084 588
rect 14140 532 14150 588
rect 11508 522 11564 532
rect 13412 522 13468 532
rect 15092 522 15148 532
rect 15204 588 15260 598
rect 16660 588 16716 598
rect 16329 537 16487 583
rect 15204 522 15260 532
rect 16660 522 16716 532
rect 17556 588 17612 598
rect 17556 522 17612 532
rect 18340 588 18396 598
rect 18340 522 18396 532
rect 18900 588 18956 598
rect 21130 532 21140 588
rect 21196 532 21206 588
rect 18900 522 18956 532
rect 14532 476 14588 486
rect 1642 420 1652 476
rect 1708 420 1718 476
rect 1866 420 1876 476
rect 1932 420 1942 476
rect 3882 420 3892 476
rect 3948 420 3958 476
rect 7354 420 7364 476
rect 7420 420 7430 476
rect 7578 420 7588 476
rect 7644 420 7654 476
rect 10154 364 10230 451
rect 12297 425 12679 471
rect 13066 420 13076 476
rect 13132 420 13142 476
rect 14313 425 14532 471
rect 14532 410 14588 420
rect 10154 308 10164 364
rect 10220 308 10230 364
rect 14746 364 14822 451
rect 15494 420 15540 476
rect 15596 420 15606 476
rect 15866 420 15876 476
rect 15932 471 15942 476
rect 18106 471 18116 476
rect 15932 425 16090 471
rect 18009 425 18116 471
rect 15932 420 15942 425
rect 18106 420 18116 425
rect 18172 420 18182 476
rect 14746 308 14756 364
rect 14812 308 14822 364
rect 18554 364 18630 451
rect 22362 420 22372 476
rect 22428 420 22438 476
rect 22586 420 22596 476
rect 22652 420 22662 476
rect 18554 308 18564 364
rect 18620 308 18630 364
rect 19338 364 19414 405
rect 19338 308 19348 364
rect 19404 308 19414 364
rect 5992 28 6044 84
rect 6100 28 6200 84
rect 6256 28 6356 84
rect 6412 28 6512 84
rect 6568 28 6668 84
rect 6724 28 6776 84
<< via1 >>
rect 16460 20636 16516 20692
rect 16616 20636 16672 20692
rect 16772 20636 16828 20692
rect 16928 20636 16984 20692
rect 17084 20636 17140 20692
rect 4116 20468 4172 20524
rect 3332 20356 3388 20412
rect 20468 20356 20524 20412
rect 2548 20244 2604 20300
rect 3668 20244 3724 20300
rect 4004 20264 4060 20320
rect 4340 20244 4396 20300
rect 4452 20244 4508 20300
rect 4676 20244 4732 20300
rect 5012 20244 5068 20300
rect 5348 20244 5404 20300
rect 6020 20244 6076 20300
rect 6356 20244 6412 20300
rect 10276 20244 10332 20300
rect 11956 20244 12012 20300
rect 12292 20244 12348 20300
rect 14084 20244 14140 20300
rect 14308 20244 14364 20300
rect 18116 20244 18172 20300
rect 19348 20244 19404 20300
rect 21140 20244 21196 20300
rect 22372 20244 22428 20300
rect 23156 20244 23212 20300
rect 1092 20132 1148 20188
rect 1316 20132 1372 20188
rect 3780 20132 3836 20188
rect 4116 20132 4172 20188
rect 8820 20132 8876 20188
rect 9044 20132 9100 20188
rect 10948 20132 11004 20188
rect 12740 20132 12796 20188
rect 13076 20132 13132 20188
rect 13636 20132 13692 20188
rect 16772 20132 16828 20188
rect 16996 20132 17052 20188
rect 18788 20132 18844 20188
rect 19908 20132 19964 20188
rect 4900 20020 4956 20076
rect 6244 20020 6300 20076
rect 22260 20132 22316 20188
rect 21476 20020 21532 20076
rect 22820 20020 22876 20076
rect 23492 20020 23548 20076
rect 12852 19908 12908 19964
rect 13300 19908 13356 19964
rect 6044 19740 6100 19796
rect 6200 19740 6256 19796
rect 6356 19740 6412 19796
rect 6512 19740 6568 19796
rect 6668 19740 6724 19796
rect 4228 19572 4284 19628
rect 21588 19572 21644 19628
rect 22820 19552 22876 19608
rect 19348 19460 19404 19516
rect 1876 19348 1932 19404
rect 1988 19348 2044 19404
rect 2996 19348 3052 19404
rect 9156 19348 9212 19404
rect 9380 19348 9436 19404
rect 11620 19348 11676 19404
rect 12628 19348 12684 19404
rect 12740 19348 12796 19404
rect 15428 19348 15484 19404
rect 15652 19348 15708 19404
rect 4116 19236 4172 19292
rect 4452 19236 4508 19292
rect 4564 19236 4620 19292
rect 4788 19256 4844 19312
rect 5348 19236 5404 19292
rect 8036 19236 8092 19292
rect 16772 19236 16828 19292
rect 18788 19236 18844 19292
rect 19124 19236 19180 19292
rect 19460 19236 19516 19292
rect 19796 19236 19852 19292
rect 21588 19236 21644 19292
rect 22820 19236 22876 19292
rect 84 19124 140 19180
rect 3892 19124 3948 19180
rect 5124 19124 5180 19180
rect 7140 19124 7196 19180
rect 11060 19124 11116 19180
rect 17444 19124 17500 19180
rect 20692 19124 20748 19180
rect 20804 19124 20860 19180
rect 22148 19124 22204 19180
rect 23604 19124 23660 19180
rect 4788 19012 4844 19068
rect 16460 18844 16516 18900
rect 16616 18844 16672 18900
rect 16772 18844 16828 18900
rect 16928 18844 16984 18900
rect 17084 18844 17140 18900
rect 420 18676 476 18732
rect 4116 18676 4172 18732
rect 84 18569 140 18625
rect 4900 18676 4956 18732
rect 7364 18676 7420 18732
rect 11844 18676 11900 18732
rect 5796 18564 5852 18620
rect 12404 18676 12460 18732
rect 15316 18676 15372 18732
rect 20356 18564 20412 18620
rect 21700 18564 21756 18620
rect 756 18452 812 18508
rect 1988 18452 2044 18508
rect 2660 18452 2716 18508
rect 3444 18452 3500 18508
rect 3668 18452 3724 18508
rect 3780 18452 3836 18508
rect 4452 18452 4508 18508
rect 4676 18452 4732 18508
rect 5124 18452 5180 18508
rect 5236 18452 5292 18508
rect 5572 18452 5628 18508
rect 5684 18452 5740 18508
rect 6132 18452 6188 18508
rect 6244 18452 6300 18508
rect 6356 18452 6412 18508
rect 6468 18452 6524 18508
rect 7588 18452 7644 18508
rect 7700 18452 7756 18508
rect 10276 18452 10332 18508
rect 11620 18452 11676 18508
rect 12740 18452 12796 18508
rect 14532 18452 14588 18508
rect 14756 18452 14812 18508
rect 15092 18452 15148 18508
rect 17332 18452 17388 18508
rect 19796 18452 19852 18508
rect 20468 18452 20524 18508
rect 21140 18452 21196 18508
rect 21812 18452 21868 18508
rect 22484 18452 22540 18508
rect 3108 18340 3164 18396
rect 4900 18340 4956 18396
rect 5908 18340 5964 18396
rect 7364 18340 7420 18396
rect 8932 18340 8988 18396
rect 9156 18340 9212 18396
rect 10948 18340 11004 18396
rect 13748 18340 13804 18396
rect 14420 18340 14476 18396
rect 16548 18340 16604 18396
rect 18452 18340 18508 18396
rect 18676 18340 18732 18396
rect 23156 18340 23212 18396
rect 196 18228 252 18284
rect 1540 18228 1596 18284
rect 4116 18228 4172 18284
rect 4564 18228 4620 18284
rect 12292 18228 12348 18284
rect 12964 18228 13020 18284
rect 20916 18228 20972 18284
rect 22260 18228 22316 18284
rect 22932 18228 22988 18284
rect 6044 17948 6100 18004
rect 6200 17948 6256 18004
rect 6356 17948 6412 18004
rect 6512 17948 6568 18004
rect 6668 17948 6724 18004
rect 19012 17668 19068 17724
rect 4228 17556 4284 17612
rect 6804 17556 6860 17612
rect 7028 17556 7084 17612
rect 11060 17556 11116 17612
rect 11284 17556 11340 17612
rect 15428 17556 15484 17612
rect 15652 17556 15708 17612
rect 420 17444 476 17500
rect 1652 17444 1708 17500
rect 2100 17444 2156 17500
rect 2548 17444 2604 17500
rect 2660 17444 2716 17500
rect 3108 17444 3164 17500
rect 3220 17444 3276 17500
rect 3556 17444 3612 17500
rect 3668 17444 3724 17500
rect 4116 17444 4172 17500
rect 8260 17444 8316 17500
rect 9380 17444 9436 17500
rect 9716 17444 9772 17500
rect 12404 17444 12460 17500
rect 16884 17444 16940 17500
rect 20244 17444 20300 17500
rect 21476 17444 21532 17500
rect 22708 17444 22764 17500
rect 196 17332 252 17388
rect 9044 17332 9100 17388
rect 9940 17332 9996 17388
rect 13300 17332 13356 17388
rect 17668 17332 17724 17388
rect 18788 17332 18844 17388
rect 19572 17332 19628 17388
rect 20804 17332 20860 17388
rect 21364 17332 21420 17388
rect 22036 17332 22092 17388
rect 22596 17332 22652 17388
rect 23716 17332 23772 17388
rect 756 17210 812 17266
rect 1876 17220 1932 17276
rect 2324 17220 2380 17276
rect 3108 17220 3164 17276
rect 3230 17220 3286 17276
rect 3892 17220 3948 17276
rect 16460 17052 16516 17108
rect 16616 17052 16672 17108
rect 16772 17052 16828 17108
rect 16928 17052 16984 17108
rect 17084 17052 17140 17108
rect 8820 16884 8876 16940
rect 9492 16884 9548 16940
rect 11060 16884 11116 16940
rect 14756 16884 14812 16940
rect 16884 16884 16940 16940
rect 4228 16772 4284 16828
rect 14644 16772 14700 16828
rect 23380 16772 23436 16828
rect 644 16660 700 16716
rect 1540 16660 1596 16716
rect 1652 16660 1708 16716
rect 1764 16660 1820 16716
rect 2100 16660 2156 16716
rect 2212 16660 2268 16716
rect 2324 16660 2380 16716
rect 2436 16660 2492 16716
rect 2548 16645 2604 16701
rect 2884 16660 2940 16716
rect 3556 16660 3612 16716
rect 3780 16660 3836 16716
rect 3892 16660 3948 16716
rect 4116 16660 4172 16716
rect 4564 16660 4620 16716
rect 5460 16660 5516 16716
rect 5908 16660 5964 16716
rect 6020 16660 6076 16716
rect 7364 16660 7420 16716
rect 7588 16660 7644 16716
rect 7700 16660 7756 16716
rect 7924 16660 7980 16716
rect 8148 16660 8204 16716
rect 8377 16660 8433 16716
rect 8489 16660 8545 16716
rect 8932 16660 8988 16716
rect 9044 16660 9100 16716
rect 9268 16660 9324 16716
rect 9716 16670 9772 16726
rect 10836 16660 10892 16716
rect 14084 16660 14140 16716
rect 14980 16660 15036 16716
rect 16660 16660 16716 16716
rect 22260 16660 22316 16716
rect 1876 16548 1932 16604
rect 5348 16548 5404 16604
rect 5796 16548 5852 16604
rect 7252 16543 7308 16599
rect 9828 16543 9884 16599
rect 10276 16548 10332 16604
rect 12740 16548 12796 16604
rect 12964 16548 13020 16604
rect 15540 16548 15596 16604
rect 16100 16548 16156 16604
rect 19348 16548 19404 16604
rect 19460 16548 19516 16604
rect 20468 16548 20524 16604
rect 21140 16548 21196 16604
rect 22148 16548 22204 16604
rect 1092 16436 1148 16492
rect 2772 16436 2828 16492
rect 6804 16436 6860 16492
rect 22708 16436 22764 16492
rect 3556 16324 3612 16380
rect 10052 16324 10108 16380
rect 15652 16324 15708 16380
rect 6044 16156 6100 16212
rect 6200 16156 6256 16212
rect 6356 16156 6412 16212
rect 6512 16156 6568 16212
rect 6668 16156 6724 16212
rect 5796 15988 5852 16044
rect 6356 15988 6412 16044
rect 13748 15988 13804 16044
rect 4340 15876 4396 15932
rect 1092 15764 1148 15820
rect 2884 15764 2940 15820
rect 3108 15764 3164 15820
rect 7812 15876 7868 15932
rect 12740 15876 12796 15932
rect 20356 15876 20412 15932
rect 9268 15764 9324 15820
rect 9492 15764 9548 15820
rect 13524 15764 13580 15820
rect 17780 15764 17836 15820
rect 18788 15764 18844 15820
rect 18900 15764 18956 15820
rect 1652 15652 1708 15708
rect 4900 15652 4956 15708
rect 5348 15652 5404 15708
rect 5572 15652 5628 15708
rect 5796 15652 5852 15708
rect 6020 15652 6076 15708
rect 6132 15652 6188 15708
rect 6356 15652 6412 15708
rect 7364 15652 7420 15708
rect 7588 15652 7644 15708
rect 10724 15652 10780 15708
rect 11956 15652 12012 15708
rect 13076 15652 13132 15708
rect 15092 15652 15148 15708
rect 20132 15652 20188 15708
rect 21252 15652 21308 15708
rect 21812 15657 21868 15713
rect 23156 15652 23212 15708
rect 4228 15540 4284 15596
rect 4564 15540 4620 15596
rect 11508 15540 11564 15596
rect 14644 15540 14700 15596
rect 17220 15540 17276 15596
rect 21140 15540 21196 15596
rect 21812 15535 21868 15591
rect 22484 15540 22540 15596
rect 23044 15540 23100 15596
rect 23716 15540 23772 15596
rect 11844 15428 11900 15484
rect 16460 15260 16516 15316
rect 16616 15260 16672 15316
rect 16772 15260 16828 15316
rect 16928 15260 16984 15316
rect 17084 15260 17140 15316
rect 756 15092 812 15148
rect 1988 15092 2044 15148
rect 4788 15092 4844 15148
rect 644 14980 700 15036
rect 3668 14980 3724 15036
rect 4452 14995 4508 15051
rect 10388 15092 10444 15148
rect 20132 15092 20188 15148
rect 21700 15092 21756 15148
rect 6468 14980 6524 15036
rect 14308 14980 14364 15036
rect 21140 14980 21196 15036
rect 22932 14985 22988 15041
rect 23604 14980 23660 15036
rect 84 14868 140 14924
rect 196 14868 252 14924
rect 1316 14868 1372 14924
rect 1428 14868 1484 14924
rect 1652 14868 1708 14924
rect 2436 14868 2492 14924
rect 2660 14868 2716 14924
rect 3220 14868 3276 14924
rect 4116 14868 4172 14924
rect 4564 14868 4620 14924
rect 7252 14868 7308 14924
rect 9940 14868 9996 14924
rect 11732 14868 11788 14924
rect 18340 14868 18396 14924
rect 22372 14868 22428 14924
rect 22932 14863 22988 14919
rect 1092 14756 1148 14812
rect 2772 14756 2828 14812
rect 4788 14756 4844 14812
rect 3780 14644 3836 14700
rect 8484 14756 8540 14812
rect 8708 14756 8764 14812
rect 10052 14756 10108 14812
rect 10500 14756 10556 14812
rect 12964 14756 13020 14812
rect 13188 14756 13244 14812
rect 16996 14756 17052 14812
rect 17220 14756 17276 14812
rect 19012 14756 19068 14812
rect 6804 14644 6860 14700
rect 11172 14644 11228 14700
rect 14532 14644 14588 14700
rect 6044 14364 6100 14420
rect 6200 14364 6256 14420
rect 6356 14364 6412 14420
rect 6512 14364 6568 14420
rect 6668 14364 6724 14420
rect 9380 14196 9436 14252
rect 3108 14089 3164 14145
rect 4228 14084 4284 14140
rect 6132 14084 6188 14140
rect 8372 14084 8428 14140
rect 16212 14084 16268 14140
rect 1092 13972 1148 14028
rect 1316 13972 1372 14028
rect 3332 13972 3388 14028
rect 3892 13972 3948 14028
rect 4900 13972 4956 14028
rect 5236 13972 5292 14028
rect 7924 13972 7980 14028
rect 12740 13972 12796 14028
rect 14532 13967 14588 14023
rect 14756 13972 14812 14028
rect 18788 13972 18844 14028
rect 18900 13972 18956 14028
rect 19908 13972 19964 14028
rect 22820 13972 22876 14028
rect 2548 13860 2604 13916
rect 3108 13860 3164 13916
rect 3668 13860 3724 13916
rect 4004 13860 4060 13916
rect 4564 13860 4620 13916
rect 4676 13860 4732 13916
rect 5796 13860 5852 13916
rect 6244 13860 6300 13916
rect 7364 13860 7420 13916
rect 7476 13860 7532 13916
rect 7700 13860 7756 13916
rect 9492 13860 9548 13916
rect 9716 13860 9772 13916
rect 10388 13860 10444 13916
rect 10612 13860 10668 13916
rect 12068 13860 12124 13916
rect 13300 13860 13356 13916
rect 15988 13880 16044 13936
rect 16436 13860 16492 13916
rect 16548 13860 16604 13916
rect 22260 13860 22316 13916
rect 2996 13748 3052 13804
rect 6020 13636 6076 13692
rect 9380 13636 9436 13692
rect 12852 13748 12908 13804
rect 17556 13748 17612 13804
rect 20804 13748 20860 13804
rect 22148 13748 22204 13804
rect 22932 13748 22988 13804
rect 10836 13636 10892 13692
rect 16460 13468 16516 13524
rect 16616 13468 16672 13524
rect 16772 13468 16828 13524
rect 16928 13468 16984 13524
rect 17084 13468 17140 13524
rect 1876 13300 1932 13356
rect 2772 13300 2828 13356
rect 3668 13300 3724 13356
rect 4228 13300 4284 13356
rect 11844 13300 11900 13356
rect 12964 13300 13020 13356
rect 19124 13300 19180 13356
rect 20580 13300 20636 13356
rect 1540 13188 1596 13244
rect 9044 13188 9100 13244
rect 18788 13188 18844 13244
rect 196 13076 252 13132
rect 1092 13076 1148 13132
rect 2212 13076 2268 13132
rect 2324 13076 2380 13132
rect 3332 13076 3388 13132
rect 3444 13076 3500 13132
rect 4116 13076 4172 13132
rect 4340 13076 4396 13132
rect 4676 13076 4732 13132
rect 8484 13076 8540 13132
rect 10500 13076 10556 13132
rect 11620 13076 11676 13132
rect 12740 13076 12796 13132
rect 14084 13076 14140 13132
rect 18116 13076 18172 13132
rect 19460 13076 19516 13132
rect 19572 13076 19628 13132
rect 20132 13076 20188 13132
rect 20244 13076 20300 13132
rect 21028 13076 21084 13132
rect 21364 13076 21420 13132
rect 22148 13076 22204 13132
rect 22932 13076 22988 13132
rect 1764 12964 1820 13020
rect 2436 12964 2492 13020
rect 7140 12964 7196 13020
rect 7364 12964 7420 13020
rect 532 12852 588 12908
rect 868 12852 924 12908
rect 4564 12852 4620 12908
rect 11172 12964 11228 13020
rect 12180 12964 12236 13020
rect 15316 12964 15372 13020
rect 15540 12964 15596 13020
rect 17556 12964 17612 13020
rect 18788 12964 18844 13020
rect 20692 12964 20748 13020
rect 21476 12969 21532 13025
rect 10052 12852 10108 12908
rect 10724 12852 10780 12908
rect 13412 12852 13468 12908
rect 18004 12852 18060 12908
rect 22596 12852 22652 12908
rect 23268 12852 23324 12908
rect 2996 12740 3052 12796
rect 9828 12740 9884 12796
rect 10836 12740 10892 12796
rect 11956 12740 12012 12796
rect 6044 12572 6100 12628
rect 6200 12572 6256 12628
rect 6356 12572 6412 12628
rect 6512 12572 6568 12628
rect 6668 12572 6724 12628
rect 4564 12404 4620 12460
rect 5572 12404 5628 12460
rect 13524 12404 13580 12460
rect 13748 12404 13804 12460
rect 14868 12404 14924 12460
rect 18228 12404 18284 12460
rect 22932 12404 22988 12460
rect 6916 12292 6972 12348
rect 8708 12292 8764 12348
rect 8820 12292 8876 12348
rect 1092 12180 1148 12236
rect 1316 12180 1372 12236
rect 3556 12180 3612 12236
rect 4452 12180 4508 12236
rect 7588 12190 7644 12246
rect 8036 12180 8092 12236
rect 8372 12180 8428 12236
rect 9604 12292 9660 12348
rect 12628 12292 12684 12348
rect 14756 12292 14812 12348
rect 16884 12292 16940 12348
rect 18004 12292 18060 12348
rect 19124 12292 19180 12348
rect 20132 12292 20188 12348
rect 11284 12180 11340 12236
rect 11508 12180 11564 12236
rect 13412 12180 13468 12236
rect 14084 12180 14140 12236
rect 15092 12180 15148 12236
rect 19796 12180 19852 12236
rect 2436 12068 2492 12124
rect 3220 12068 3276 12124
rect 3892 12068 3948 12124
rect 5684 12068 5740 12124
rect 5796 12068 5852 12124
rect 7476 12068 7532 12124
rect 7812 12078 7868 12134
rect 8596 12068 8652 12124
rect 9044 12068 9100 12124
rect 9156 12068 9212 12124
rect 10164 12068 10220 12124
rect 12964 12068 13020 12124
rect 14420 12068 14476 12124
rect 15540 12068 15596 12124
rect 15876 12068 15932 12124
rect 17556 12088 17612 12144
rect 18564 12068 18620 12124
rect 19236 12068 19292 12124
rect 20468 12068 20524 12124
rect 20692 12068 20748 12124
rect 21700 12068 21756 12124
rect 21924 12068 21980 12124
rect 22596 12063 22652 12119
rect 5348 11956 5404 12012
rect 7700 11956 7756 12012
rect 7924 11951 7980 12007
rect 19796 11956 19852 12012
rect 21476 11956 21532 12012
rect 22820 11956 22876 12012
rect 6244 11844 6300 11900
rect 16460 11676 16516 11732
rect 16616 11676 16672 11732
rect 16772 11676 16828 11732
rect 16928 11676 16984 11732
rect 17084 11676 17140 11732
rect 5236 11396 5292 11452
rect 21252 11396 21308 11452
rect 22148 11401 22204 11457
rect 2996 11284 3052 11340
rect 4004 11284 4060 11340
rect 4340 11284 4396 11340
rect 4676 11284 4732 11340
rect 7700 11284 7756 11340
rect 12852 11284 12908 11340
rect 13748 11284 13804 11340
rect 17108 11284 17164 11340
rect 20244 11284 20300 11340
rect 21588 11284 21644 11340
rect 22148 11279 22204 11335
rect 1652 11172 1708 11228
rect 1876 11172 1932 11228
rect 3780 11172 3836 11228
rect 4564 11172 4620 11228
rect 6916 11172 6972 11228
rect 8932 11172 8988 11228
rect 9156 11172 9212 11228
rect 11508 11172 11564 11228
rect 11732 11172 11788 11228
rect 13412 11172 13468 11228
rect 14196 11172 14252 11228
rect 16212 11172 16268 11228
rect 18228 11172 18284 11228
rect 18452 11172 18508 11228
rect 20020 11172 20076 11228
rect 20804 11172 20860 11228
rect 22820 11172 22876 11228
rect 5236 11060 5292 11116
rect 13524 11060 13580 11116
rect 19908 11060 19964 11116
rect 21028 11060 21084 11116
rect 23268 11060 23324 11116
rect 14420 10948 14476 11004
rect 6044 10780 6100 10836
rect 6200 10780 6256 10836
rect 6356 10780 6412 10836
rect 6512 10780 6568 10836
rect 6668 10780 6724 10836
rect 12740 10612 12796 10668
rect 13412 10612 13468 10668
rect 532 10500 588 10556
rect 11732 10500 11788 10556
rect 14532 10500 14588 10556
rect 15428 10500 15484 10556
rect 17444 10500 17500 10556
rect 18676 10500 18732 10556
rect 756 10388 812 10444
rect 2752 10388 2808 10444
rect 2996 10388 3052 10444
rect 4116 10388 4172 10444
rect 6020 10388 6076 10444
rect 6244 10388 6300 10444
rect 9716 10388 9772 10444
rect 9940 10388 9996 10444
rect 11620 10388 11676 10444
rect 12404 10388 12460 10444
rect 13636 10388 13692 10444
rect 14308 10388 14364 10444
rect 14868 10388 14924 10444
rect 15876 10388 15932 10444
rect 16212 10388 16268 10444
rect 196 10276 252 10332
rect 980 10276 1036 10332
rect 1204 10276 1260 10332
rect 1428 10276 1484 10332
rect 1652 10276 1708 10332
rect 2324 10276 2380 10332
rect 3220 10276 3276 10332
rect 3332 10276 3388 10332
rect 4788 10276 4844 10332
rect 11060 10276 11116 10332
rect 11956 10276 12012 10332
rect 3556 10164 3612 10220
rect 14196 10276 14252 10332
rect 15092 10276 15148 10332
rect 15428 10276 15484 10332
rect 18340 10383 18396 10439
rect 20020 10388 20076 10444
rect 20468 10388 20524 10444
rect 22372 10388 22428 10444
rect 22596 10388 22652 10444
rect 15988 10276 16044 10332
rect 16324 10276 16380 10332
rect 18228 10276 18284 10332
rect 19348 10296 19404 10352
rect 19460 10276 19516 10332
rect 21140 10276 21196 10332
rect 3668 10164 3724 10220
rect 19796 10164 19852 10220
rect 1652 10052 1708 10108
rect 15204 10052 15260 10108
rect 16460 9884 16516 9940
rect 16616 9884 16672 9940
rect 16772 9884 16828 9940
rect 16928 9884 16984 9940
rect 17084 9884 17140 9940
rect 644 9716 700 9772
rect 980 9716 1036 9772
rect 1316 9716 1372 9772
rect 11732 9716 11788 9772
rect 11844 9716 11900 9772
rect 14756 9716 14812 9772
rect 14980 9716 15036 9772
rect 22484 9716 22540 9772
rect 10164 9604 10220 9660
rect 15988 9604 16044 9660
rect 23716 9604 23772 9660
rect 84 9492 140 9548
rect 756 9497 812 9553
rect 1204 9492 1260 9548
rect 1540 9482 1596 9538
rect 1876 9492 1932 9548
rect 1988 9492 2044 9548
rect 2660 9487 2716 9543
rect 3892 9497 3948 9553
rect 4116 9492 4172 9548
rect 4676 9492 4732 9548
rect 7924 9492 7980 9548
rect 9268 9492 9324 9548
rect 9828 9492 9884 9548
rect 10612 9492 10668 9548
rect 11508 9492 11564 9548
rect 12180 9492 12236 9548
rect 12964 9492 13020 9548
rect 13748 9492 13804 9548
rect 13972 9492 14028 9548
rect 14084 9492 14140 9548
rect 14196 9492 14252 9548
rect 14532 9492 14588 9548
rect 14644 9492 14700 9548
rect 14868 9497 14924 9553
rect 14980 9492 15036 9548
rect 15540 9502 15596 9558
rect 15652 9492 15708 9548
rect 17108 9492 17164 9548
rect 19684 9492 19740 9548
rect 22260 9492 22316 9548
rect 22932 9492 22988 9548
rect 644 9370 700 9426
rect 2660 9365 2716 9421
rect 3444 9380 3500 9436
rect 3668 9380 3724 9436
rect 3780 9355 3836 9411
rect 4228 9360 4284 9416
rect 6580 9380 6636 9436
rect 6804 9380 6860 9436
rect 8596 9380 8652 9436
rect 9940 9380 9996 9436
rect 10948 9380 11004 9436
rect 12628 9380 12684 9436
rect 16100 9380 16156 9436
rect 17668 9380 17724 9436
rect 2324 9268 2380 9324
rect 17892 9380 17948 9436
rect 18788 9380 18844 9436
rect 20804 9380 20860 9436
rect 21028 9380 21084 9436
rect 15540 9268 15596 9324
rect 17332 9268 17388 9324
rect 10724 9156 10780 9212
rect 12740 9156 12796 9212
rect 6044 8988 6100 9044
rect 6200 8988 6256 9044
rect 6356 8988 6412 9044
rect 6512 8988 6568 9044
rect 6668 8988 6724 9044
rect 1204 8820 1260 8876
rect 15428 8820 15484 8876
rect 2884 8708 2940 8764
rect 5684 8708 5740 8764
rect 7028 8708 7084 8764
rect 13636 8708 13692 8764
rect 15316 8708 15372 8764
rect 16100 8708 16156 8764
rect 16324 8708 16380 8764
rect 16772 8708 16828 8764
rect 17546 8708 17602 8764
rect 17892 8708 17948 8764
rect 19236 8708 19292 8764
rect 308 8596 364 8652
rect 980 8596 1036 8652
rect 2436 8596 2492 8652
rect 2996 8596 3052 8652
rect 3556 8596 3612 8652
rect 9604 8596 9660 8652
rect 11060 8596 11116 8652
rect 11284 8596 11340 8652
rect 13300 8596 13356 8652
rect 17780 8596 17836 8652
rect 19572 8708 19628 8764
rect 20132 8708 20188 8764
rect 23492 8713 23548 8769
rect 20580 8596 20636 8652
rect 1092 8484 1148 8540
rect 2660 8484 2716 8540
rect 2772 8484 2828 8540
rect 3108 8484 3164 8540
rect 3332 8484 3388 8540
rect 3780 8484 3836 8540
rect 3892 8484 3948 8540
rect 4116 8494 4172 8550
rect 84 8372 140 8428
rect 3444 8372 3500 8428
rect 4340 8427 4396 8483
rect 5460 8484 5516 8540
rect 5572 8484 5628 8540
rect 5796 8484 5852 8540
rect 5908 8484 5964 8540
rect 6916 8484 6972 8540
rect 7252 8484 7308 8540
rect 7364 8484 7420 8540
rect 7700 8484 7756 8540
rect 8036 8484 8092 8540
rect 8148 8484 8204 8540
rect 9268 8464 9324 8520
rect 9380 8484 9436 8540
rect 12516 8484 12572 8540
rect 14420 8484 14476 8540
rect 14644 8484 14700 8540
rect 14756 8484 14812 8540
rect 15204 8484 15260 8540
rect 15428 8484 15484 8540
rect 15652 8489 15708 8545
rect 15764 8484 15820 8540
rect 18228 8484 18284 8540
rect 18340 8484 18396 8540
rect 18676 8484 18732 8540
rect 19684 8484 19740 8540
rect 20916 8484 20972 8540
rect 23044 8484 23100 8540
rect 5124 8372 5180 8428
rect 7476 8372 7532 8428
rect 14868 8372 14924 8428
rect 16324 8372 16380 8428
rect 17220 8372 17276 8428
rect 3556 8260 3612 8316
rect 4116 8260 4172 8316
rect 5460 8260 5516 8316
rect 7252 8260 7308 8316
rect 9716 8260 9772 8316
rect 19124 8372 19180 8428
rect 22372 8372 22428 8428
rect 18900 8260 18956 8316
rect 20692 8260 20748 8316
rect 21476 8260 21532 8316
rect 16460 8092 16516 8148
rect 16616 8092 16672 8148
rect 16772 8092 16828 8148
rect 16928 8092 16984 8148
rect 17084 8092 17140 8148
rect 5572 7924 5628 7980
rect 9380 7924 9436 7980
rect 14420 7924 14476 7980
rect 14756 7924 14812 7980
rect 15652 7924 15708 7980
rect 16212 7924 16268 7980
rect 17668 7812 17724 7868
rect 19124 7812 19180 7868
rect 19684 7812 19740 7868
rect 21140 7812 21196 7868
rect 22148 7812 22204 7868
rect 3220 7700 3276 7756
rect 4004 7700 4060 7756
rect 4452 7700 4508 7756
rect 4676 7700 4732 7756
rect 4788 7700 4844 7756
rect 5124 7700 5180 7756
rect 5796 7700 5852 7756
rect 5908 7700 5964 7756
rect 6916 7705 6972 7761
rect 7364 7700 7420 7756
rect 7608 7700 7664 7756
rect 9044 7700 9100 7756
rect 9156 7700 9212 7756
rect 9492 7700 9548 7756
rect 13076 7700 13132 7756
rect 14532 7700 14588 7756
rect 14980 7700 15036 7756
rect 15876 7680 15932 7736
rect 15988 7700 16044 7756
rect 16212 7700 16268 7756
rect 16548 7700 16604 7756
rect 17780 7700 17836 7756
rect 18228 7700 18284 7756
rect 18340 7700 18396 7756
rect 19908 7700 19964 7756
rect 21364 7700 21420 7756
rect 21476 7700 21532 7756
rect 1876 7588 1932 7644
rect 2100 7588 2156 7644
rect 6916 7583 6972 7639
rect 10052 7588 10108 7644
rect 11732 7588 11788 7644
rect 11956 7588 12012 7644
rect 15652 7588 15708 7644
rect 16100 7588 16156 7644
rect 22708 7700 22764 7756
rect 17444 7588 17500 7644
rect 18004 7588 18060 7644
rect 8260 7476 8316 7532
rect 8708 7476 8764 7532
rect 13636 7476 13692 7532
rect 18676 7476 18732 7532
rect 19348 7588 19404 7644
rect 20916 7588 20972 7644
rect 22148 7588 22204 7644
rect 23380 7588 23436 7644
rect 19572 7476 19628 7532
rect 21812 7476 21868 7532
rect 22932 7476 22988 7532
rect 7364 7364 7420 7420
rect 17444 7364 17500 7420
rect 18004 7364 18060 7420
rect 6044 7196 6100 7252
rect 6200 7196 6256 7252
rect 6356 7196 6412 7252
rect 6512 7196 6568 7252
rect 6668 7196 6724 7252
rect 13188 7028 13244 7084
rect 14756 7028 14812 7084
rect 12740 6916 12796 6972
rect 15652 6916 15708 6972
rect 17780 6936 17836 6992
rect 1876 6804 1932 6860
rect 2100 6804 2156 6860
rect 3892 6804 3948 6860
rect 5796 6804 5852 6860
rect 6132 6804 6188 6860
rect 7700 6804 7756 6860
rect 8596 6804 8652 6860
rect 10612 6804 10668 6860
rect 10836 6804 10892 6860
rect 12516 6814 12572 6870
rect 13300 6804 13356 6860
rect 13972 6804 14028 6860
rect 14756 6804 14812 6860
rect 16212 6819 16268 6875
rect 18004 6814 18060 6870
rect 19012 6824 19068 6880
rect 19124 6809 19180 6865
rect 22036 6804 22092 6860
rect 3220 6692 3276 6748
rect 4676 6692 4732 6748
rect 5124 6692 5180 6748
rect 5236 6692 5292 6748
rect 5460 6692 5516 6748
rect 5684 6692 5740 6748
rect 7812 6692 7868 6748
rect 8260 6692 8316 6748
rect 9492 6692 9548 6748
rect 11956 6687 12012 6743
rect 12628 6692 12684 6748
rect 12964 6692 13020 6748
rect 13860 6692 13916 6748
rect 14980 6692 15036 6748
rect 15092 6692 15148 6748
rect 15540 6692 15596 6748
rect 15764 6692 15820 6748
rect 16324 6697 16380 6753
rect 17668 6692 17724 6748
rect 17892 6692 17948 6748
rect 19348 6692 19404 6748
rect 19684 6692 19740 6748
rect 19908 6692 19964 6748
rect 15988 6580 16044 6636
rect 16660 6580 16716 6636
rect 20356 6692 20412 6748
rect 20468 6692 20524 6748
rect 20692 6692 20748 6748
rect 21028 6692 21084 6748
rect 21588 6692 21644 6748
rect 22820 6692 22876 6748
rect 23716 6692 23772 6748
rect 18228 6580 18284 6636
rect 19236 6580 19292 6636
rect 19460 6580 19516 6636
rect 3780 6468 3836 6524
rect 4564 6468 4620 6524
rect 4900 6468 4956 6524
rect 8036 6468 8092 6524
rect 12516 6468 12572 6524
rect 16324 6458 16380 6514
rect 20020 6468 20076 6524
rect 21252 6468 21308 6524
rect 21924 6468 21980 6524
rect 16460 6300 16516 6356
rect 16616 6300 16672 6356
rect 16772 6300 16828 6356
rect 16928 6300 16984 6356
rect 17084 6300 17140 6356
rect 4228 6132 4284 6188
rect 4798 6132 4854 6188
rect 5572 6132 5628 6188
rect 6020 6132 6076 6188
rect 6916 6132 6972 6188
rect 7476 6132 7532 6188
rect 3892 6020 3948 6076
rect 5236 6020 5292 6076
rect 8036 6020 8092 6076
rect 14186 6030 14242 6086
rect 14532 6020 14588 6076
rect 16660 6020 16716 6076
rect 18564 6020 18620 6076
rect 20356 6015 20412 6071
rect 3108 5908 3164 5964
rect 4452 5908 4508 5964
rect 4564 5903 4620 5959
rect 5012 5908 5068 5964
rect 5348 5908 5404 5964
rect 5796 5908 5852 5964
rect 6916 5908 6972 5964
rect 7140 5908 7196 5964
rect 7252 5908 7308 5964
rect 7588 5908 7644 5964
rect 10500 5908 10556 5964
rect 12404 5908 12460 5964
rect 12516 5913 12572 5969
rect 13636 5908 13692 5964
rect 14196 5903 14252 5959
rect 14644 5908 14700 5964
rect 16100 5908 16156 5964
rect 17556 5908 17612 5964
rect 19236 5908 19292 5964
rect 19348 5908 19404 5964
rect 1652 5796 1708 5852
rect 1876 5796 1932 5852
rect 9156 5796 9212 5852
rect 9380 5796 9436 5852
rect 11284 5796 11340 5852
rect 12740 5801 12796 5857
rect 12964 5796 13020 5852
rect 15428 5796 15484 5852
rect 18340 5796 18396 5852
rect 21252 5796 21308 5852
rect 22260 5796 22316 5852
rect 22372 5796 22428 5852
rect 7364 5684 7420 5740
rect 12628 5679 12684 5735
rect 13524 5684 13580 5740
rect 15876 5684 15932 5740
rect 18004 5684 18060 5740
rect 18900 5659 18956 5715
rect 6044 5404 6100 5460
rect 6200 5404 6256 5460
rect 6356 5404 6412 5460
rect 6512 5404 6568 5460
rect 6668 5404 6724 5460
rect 9716 5241 9772 5297
rect 11396 5236 11452 5292
rect 12628 5236 12684 5292
rect 2324 5124 2380 5180
rect 5124 5124 5180 5180
rect 10164 5124 10220 5180
rect 12740 5124 12796 5180
rect 17780 5124 17836 5180
rect 2884 5012 2940 5068
rect 3220 5012 3276 5068
rect 4004 5012 4060 5068
rect 4116 5012 4172 5068
rect 4564 5012 4620 5068
rect 4676 5022 4732 5078
rect 4900 5012 4956 5068
rect 9604 4992 9660 5048
rect 11284 5012 11340 5068
rect 12404 5012 12460 5068
rect 14644 5012 14700 5068
rect 15652 5030 15708 5086
rect 17220 5012 17276 5068
rect 18676 5012 18732 5068
rect 19012 5012 19068 5068
rect 20356 5012 20412 5068
rect 20580 5012 20636 5068
rect 22484 5012 22540 5068
rect 84 4900 140 4956
rect 420 4900 476 4956
rect 1092 4900 1148 4956
rect 1540 4900 1596 4956
rect 1764 4900 1820 4956
rect 1876 4900 1932 4956
rect 2100 4900 2156 4956
rect 2212 4900 2268 4956
rect 2436 4900 2492 4956
rect 2660 4900 2716 4956
rect 2996 4900 3052 4956
rect 3332 4900 3388 4956
rect 3444 4900 3500 4956
rect 3892 4900 3948 4956
rect 5460 4900 5516 4956
rect 5572 4900 5628 4956
rect 5684 4900 5740 4956
rect 6132 4900 6188 4956
rect 6356 4900 6412 4956
rect 7252 4900 7308 4956
rect 8036 4900 8092 4956
rect 8372 4900 8428 4956
rect 8484 4900 8540 4956
rect 8596 4900 8652 4956
rect 9156 4900 9212 4956
rect 10836 4900 10892 4956
rect 11956 4900 12012 4956
rect 12964 4900 13020 4956
rect 13412 4905 13468 4961
rect 13636 4900 13692 4956
rect 13860 4900 13916 4956
rect 13972 4900 14028 4956
rect 14868 4900 14924 4956
rect 15311 4900 15367 4956
rect 15540 4890 15596 4946
rect 15764 4900 15820 4956
rect 17556 4900 17612 4956
rect 18116 4900 18172 4956
rect 21700 4900 21756 4956
rect 22932 4900 22988 4956
rect 23716 4900 23772 4956
rect 5236 4788 5292 4844
rect 5908 4788 5964 4844
rect 6244 4788 6300 4844
rect 7476 4788 7532 4844
rect 14308 4788 14364 4844
rect 84 4676 140 4732
rect 2548 4676 2604 4732
rect 3668 4676 3724 4732
rect 8820 4676 8876 4732
rect 11620 4676 11676 4732
rect 18452 4676 18508 4732
rect 18788 4676 18844 4732
rect 16460 4508 16516 4564
rect 16616 4508 16672 4564
rect 16772 4508 16828 4564
rect 16928 4508 16984 4564
rect 17084 4508 17140 4564
rect 868 4340 924 4396
rect 2884 4340 2940 4396
rect 4116 4345 4172 4401
rect 4452 4340 4508 4396
rect 13412 4340 13468 4396
rect 15428 4340 15484 4396
rect 308 4228 364 4284
rect 2436 4228 2492 4284
rect 4788 4228 4844 4284
rect 17892 4228 17948 4284
rect 23492 4228 23548 4284
rect 84 4116 140 4172
rect 420 4116 476 4172
rect 980 4116 1036 4172
rect 1316 4116 1372 4172
rect 1540 4116 1596 4172
rect 1652 4116 1708 4172
rect 1876 4116 1932 4172
rect 1988 4116 2044 4172
rect 2324 4116 2380 4172
rect 2660 4116 2716 4172
rect 3108 4116 3164 4172
rect 3780 4116 3836 4172
rect 4116 4116 4172 4172
rect 4340 4116 4396 4172
rect 4564 4116 4620 4172
rect 4900 4116 4956 4172
rect 8708 4116 8764 4172
rect 12852 4116 12908 4172
rect 14308 4116 14364 4172
rect 14868 4116 14924 4172
rect 16996 4116 17052 4172
rect 17444 4116 17500 4172
rect 18340 4116 18396 4172
rect 18788 4116 18844 4172
rect 22148 4116 22204 4172
rect 23044 4116 23100 4172
rect 2212 4004 2268 4060
rect 7364 4004 7420 4060
rect 7588 4004 7644 4060
rect 9604 4004 9660 4060
rect 11508 4004 11564 4060
rect 11732 4004 11788 4060
rect 14420 4004 14476 4060
rect 15204 4004 15260 4060
rect 17892 4004 17948 4060
rect 19908 4004 19964 4060
rect 20020 4004 20076 4060
rect 21028 4004 21084 4060
rect 21588 4004 21644 4060
rect 22820 4004 22876 4060
rect 14756 3892 14812 3948
rect 17220 3892 17276 3948
rect 18564 3892 18620 3948
rect 17780 3780 17836 3836
rect 6044 3612 6100 3668
rect 6200 3612 6256 3668
rect 6356 3612 6412 3668
rect 6512 3612 6568 3668
rect 6668 3612 6724 3668
rect 4564 3444 4620 3500
rect 5012 3444 5068 3500
rect 13636 3444 13692 3500
rect 1428 3332 1484 3388
rect 4452 3337 4508 3393
rect 5796 3332 5852 3388
rect 13300 3332 13356 3388
rect 868 3220 924 3276
rect 1540 3220 1596 3276
rect 2212 3220 2268 3276
rect 3444 3220 3500 3276
rect 8260 3220 8316 3276
rect 10052 3215 10108 3271
rect 10276 3220 10332 3276
rect 12516 3220 12572 3276
rect 13860 3332 13916 3388
rect 15316 3332 15372 3388
rect 15988 3332 16044 3388
rect 17220 3332 17276 3388
rect 20244 3332 20300 3388
rect 23044 3332 23100 3388
rect 15092 3220 15148 3276
rect 17444 3220 17500 3276
rect 17780 3220 17836 3276
rect 18564 3220 18620 3276
rect 19012 3220 19068 3276
rect 20804 3220 20860 3276
rect 21476 3220 21532 3276
rect 21588 3220 21644 3276
rect 21924 3220 21980 3276
rect 23380 3220 23436 3276
rect 2436 3108 2492 3164
rect 2548 3108 2604 3164
rect 2772 3108 2828 3164
rect 3780 3108 3836 3164
rect 3892 3108 3948 3164
rect 4116 3108 4172 3164
rect 4228 3108 4284 3164
rect 4564 3108 4620 3164
rect 5236 3108 5292 3164
rect 5460 3108 5516 3164
rect 7364 3108 7420 3164
rect 7700 3108 7756 3164
rect 7924 3108 7980 3164
rect 8036 3108 8092 3164
rect 8708 3108 8764 3164
rect 8820 3108 8876 3164
rect 11508 3108 11564 3164
rect 12964 3108 13020 3164
rect 14084 3108 14140 3164
rect 14756 3103 14812 3159
rect 15316 3108 15372 3164
rect 15652 3108 15708 3164
rect 16100 3108 16156 3164
rect 16996 3108 17052 3164
rect 18116 3108 18172 3164
rect 18228 3108 18284 3164
rect 19348 3108 19404 3164
rect 20020 3108 20076 3164
rect 22484 3108 22540 3164
rect 22596 3108 22652 3164
rect 644 2996 700 3052
rect 8596 2996 8652 3052
rect 12292 2996 12348 3052
rect 14644 2996 14700 3052
rect 1876 2884 1932 2940
rect 4788 2884 4844 2940
rect 7700 2884 7756 2940
rect 8260 2884 8316 2940
rect 18788 2884 18844 2940
rect 20580 2884 20636 2940
rect 22148 2884 22204 2940
rect 16460 2716 16516 2772
rect 16616 2716 16672 2772
rect 16772 2716 16828 2772
rect 16928 2716 16984 2772
rect 17084 2716 17140 2772
rect 4228 2548 4284 2604
rect 7476 2548 7532 2604
rect 3892 2436 3948 2492
rect 5124 2436 5180 2492
rect 9268 2548 9324 2604
rect 9940 2548 9996 2604
rect 15652 2548 15708 2604
rect 18228 2548 18284 2604
rect 18676 2548 18732 2604
rect 10388 2436 10444 2492
rect 18004 2436 18060 2492
rect 3108 2324 3164 2380
rect 4452 2324 4508 2380
rect 1652 2212 1708 2268
rect 1876 2212 1932 2268
rect 5572 2324 5628 2380
rect 7700 2319 7756 2375
rect 8596 2324 8652 2380
rect 8708 2324 8764 2380
rect 8932 2324 8988 2380
rect 9156 2324 9212 2380
rect 9268 2324 9324 2380
rect 9604 2324 9660 2380
rect 9716 2324 9772 2380
rect 10164 2324 10220 2380
rect 10500 2324 10556 2380
rect 10836 2324 10892 2380
rect 11060 2324 11116 2380
rect 11732 2324 11788 2380
rect 12292 2324 12348 2380
rect 13188 2324 13244 2380
rect 13524 2324 13580 2380
rect 14196 2324 14252 2380
rect 14532 2324 14588 2380
rect 14644 2324 14700 2380
rect 14858 2324 14914 2380
rect 14980 2324 15036 2380
rect 15316 2324 15372 2380
rect 15876 2324 15932 2380
rect 15988 2324 16044 2380
rect 16212 2324 16268 2380
rect 16436 2324 16492 2380
rect 16548 2324 16604 2380
rect 16772 2324 16828 2380
rect 18116 2324 18172 2380
rect 18340 2324 18396 2380
rect 18452 2324 18508 2380
rect 18788 2324 18844 2380
rect 21028 2324 21084 2380
rect 21140 2324 21196 2380
rect 5124 2212 5180 2268
rect 6244 2212 6300 2268
rect 3668 2100 3724 2156
rect 8036 2202 8092 2258
rect 11172 2212 11228 2268
rect 14420 2212 14476 2268
rect 17668 2212 17724 2268
rect 4676 2100 4732 2156
rect 5348 2100 5404 2156
rect 8260 2095 8316 2151
rect 10612 2100 10668 2156
rect 20356 2212 20412 2268
rect 22260 2212 22316 2268
rect 22484 2212 22540 2268
rect 13524 2090 13580 2146
rect 15204 2100 15260 2156
rect 15652 2100 15708 2156
rect 19124 2100 19180 2156
rect 16772 1988 16828 2044
rect 6044 1820 6100 1876
rect 6200 1820 6256 1876
rect 6356 1820 6412 1876
rect 6512 1820 6568 1876
rect 6668 1820 6724 1876
rect 17556 1652 17612 1708
rect 2324 1540 2380 1596
rect 3556 1540 3612 1596
rect 4228 1540 4284 1596
rect 5124 1540 5180 1596
rect 5572 1540 5628 1596
rect 7700 1540 7756 1596
rect 9940 1540 9996 1596
rect 13300 1540 13356 1596
rect 13972 1540 14028 1596
rect 14532 1540 14588 1596
rect 14756 1540 14812 1596
rect 17108 1540 17164 1596
rect 308 1428 364 1484
rect 868 1428 924 1484
rect 1204 1428 1260 1484
rect 1764 1428 1820 1484
rect 2436 1428 2492 1484
rect 2996 1428 3052 1484
rect 3668 1428 3724 1484
rect 7588 1428 7644 1484
rect 15316 1428 15372 1484
rect 16212 1423 16268 1479
rect 16324 1423 16380 1479
rect 17892 1428 17948 1484
rect 18564 1428 18620 1484
rect 20244 1428 20300 1484
rect 20468 1428 20524 1484
rect 22260 1428 22316 1484
rect 196 1316 252 1372
rect 2772 1316 2828 1372
rect 4004 1316 4060 1372
rect 4340 1316 4396 1372
rect 5012 1316 5068 1372
rect 5684 1316 5740 1372
rect 6020 1316 6076 1372
rect 6356 1316 6412 1372
rect 8148 1316 8204 1372
rect 9828 1316 9884 1372
rect 10388 1316 10444 1372
rect 11396 1316 11452 1372
rect 12068 1316 12124 1372
rect 12292 1316 12348 1372
rect 12740 1316 12796 1372
rect 13076 1316 13132 1372
rect 13412 1311 13468 1367
rect 13748 1316 13804 1372
rect 14532 1316 14588 1372
rect 14980 1316 15036 1372
rect 15092 1316 15148 1372
rect 15988 1311 16044 1367
rect 18228 1316 18284 1372
rect 21588 1316 21644 1372
rect 23716 1316 23772 1372
rect 8708 1204 8764 1260
rect 12628 1204 12684 1260
rect 16460 924 16516 980
rect 16616 924 16672 980
rect 16772 924 16828 980
rect 16928 924 16984 980
rect 17084 924 17140 980
rect 4452 756 4508 812
rect 12180 756 12236 812
rect 15764 756 15820 812
rect 9268 644 9324 700
rect 20692 644 20748 700
rect 3108 532 3164 588
rect 4676 532 4732 588
rect 4900 532 4956 588
rect 8708 532 8764 588
rect 10500 532 10556 588
rect 11508 532 11564 588
rect 12852 532 12908 588
rect 13412 532 13468 588
rect 13524 532 13580 588
rect 14084 532 14140 588
rect 15092 532 15148 588
rect 15204 532 15260 588
rect 16660 532 16716 588
rect 17556 532 17612 588
rect 18340 532 18396 588
rect 18900 532 18956 588
rect 21140 532 21196 588
rect 1652 420 1708 476
rect 1876 420 1932 476
rect 3892 420 3948 476
rect 7364 420 7420 476
rect 7588 420 7644 476
rect 13076 420 13132 476
rect 14532 420 14588 476
rect 10164 308 10220 364
rect 15540 420 15596 476
rect 15876 420 15932 476
rect 18116 420 18172 476
rect 14756 308 14812 364
rect 22372 420 22428 476
rect 22596 420 22652 476
rect 18564 308 18620 364
rect 19348 308 19404 364
rect 6044 28 6100 84
rect 6200 28 6256 84
rect 6356 28 6412 84
rect 6512 28 6568 84
rect 6668 28 6724 84
<< metal2 >>
rect 4116 20524 4172 20534
rect 3332 20412 3388 20422
rect 2548 20300 2604 20310
rect 1092 20188 1148 20198
rect 1316 20188 1372 20198
rect 1148 20132 1260 20188
rect 2548 20132 2604 20244
rect 2996 20300 3052 20310
rect 1092 20122 1148 20132
rect 868 19404 924 19414
rect 84 19180 140 19190
rect 84 18625 140 19124
rect 420 18732 476 18742
rect 74 18569 84 18625
rect 140 18569 150 18625
rect 84 18503 140 18513
rect 84 14924 140 18447
rect 196 18284 252 18294
rect 196 18060 252 18228
rect 196 17994 252 18004
rect 420 17500 476 18676
rect 196 17388 252 17398
rect 196 17220 252 17332
rect 84 14858 140 14868
rect 196 14924 252 14934
rect 196 13132 252 14868
rect 196 12908 252 13076
rect 196 12842 252 12852
rect 196 10332 252 10342
rect 196 9996 252 10276
rect 196 9930 252 9940
rect 308 10108 364 10118
rect 84 9548 140 9558
rect 140 9492 252 9548
rect 84 9482 140 9492
rect 308 8652 364 10052
rect 420 9996 476 17444
rect 756 18732 812 18742
rect 756 18508 812 18676
rect 644 17388 700 17398
rect 756 17388 812 18452
rect 700 17332 812 17388
rect 644 16716 700 17332
rect 644 16650 700 16660
rect 756 17266 812 17276
rect 756 15708 812 17210
rect 756 15642 812 15652
rect 644 15596 700 15606
rect 868 15586 924 19348
rect 1316 19292 1372 20132
rect 1876 19404 1932 19414
rect 1876 19236 1932 19348
rect 1988 19404 2044 19414
rect 1988 19292 2044 19348
rect 1092 16492 1148 16502
rect 1092 16049 1148 16436
rect 1082 15993 1092 16049
rect 1148 15993 1158 16049
rect 1092 15927 1148 15937
rect 1092 15820 1148 15871
rect 1092 15754 1148 15764
rect 644 15036 700 15540
rect 756 15530 924 15586
rect 1316 15596 1372 19236
rect 1988 19226 2044 19236
rect 2996 19404 3052 20244
rect 1988 18732 2044 18742
rect 1988 18508 2044 18676
rect 1988 18442 2044 18452
rect 2660 18508 2716 18518
rect 1540 18284 1596 18294
rect 1540 17612 1596 18228
rect 1540 17546 1596 17556
rect 1652 18284 1708 18294
rect 1652 17500 1708 18228
rect 2660 17846 2716 18452
rect 2548 17790 2716 17846
rect 1540 17164 1596 17174
rect 1540 16716 1596 17108
rect 1652 17052 1708 17444
rect 2100 17500 2156 17510
rect 2548 17500 2604 17790
rect 2156 17444 2268 17500
rect 2100 17434 2156 17444
rect 1876 17276 1932 17286
rect 1876 17169 1932 17220
rect 2324 17276 2380 17286
rect 1866 17113 1876 17169
rect 1932 17113 1942 17169
rect 1866 16996 1876 17052
rect 1932 16996 1942 17052
rect 1652 16986 1708 16996
rect 1540 16650 1596 16660
rect 1652 16828 1708 16838
rect 1652 16716 1708 16772
rect 1652 15932 1708 16660
rect 1764 16716 1820 16828
rect 1764 16650 1820 16660
rect 1652 15866 1708 15876
rect 1876 16604 1932 16996
rect 2324 16940 2380 17220
rect 2324 16884 2492 16940
rect 2100 16716 2156 16726
rect 1988 16660 2100 16716
rect 2100 16650 2156 16660
rect 2212 16716 2268 16726
rect 1652 15708 1708 15805
rect 1652 15642 1708 15652
rect 1316 15530 1372 15540
rect 756 15148 812 15530
rect 756 15082 812 15092
rect 868 15464 924 15474
rect 644 14970 700 14980
rect 532 12908 588 12918
rect 532 12348 588 12852
rect 868 12908 924 15408
rect 1316 14924 1372 14934
rect 1092 14812 1148 14822
rect 1092 14160 1148 14756
rect 1316 14812 1372 14868
rect 1428 14924 1484 15036
rect 1428 14858 1484 14868
rect 1652 14924 1708 14934
rect 1316 14746 1372 14756
rect 1540 14364 1596 14374
rect 1092 14104 1260 14160
rect 1092 14028 1148 14038
rect 1092 13804 1148 13972
rect 1092 13738 1148 13748
rect 1092 13132 1148 13142
rect 1092 13020 1148 13076
rect 1092 12954 1148 12964
rect 532 12282 588 12292
rect 756 12348 812 12358
rect 532 11340 588 11350
rect 532 10556 588 11284
rect 532 10490 588 10500
rect 756 10444 812 12292
rect 756 10378 812 10388
rect 420 9930 476 9940
rect 868 9884 924 12852
rect 1204 12796 1260 14104
rect 1204 12730 1260 12740
rect 1316 14028 1372 14038
rect 1316 12348 1372 13972
rect 1092 12236 1148 12246
rect 1316 12236 1372 12292
rect 1148 12180 1260 12236
rect 1092 12170 1148 12180
rect 1316 12170 1372 12180
rect 1428 13916 1484 13926
rect 1204 11452 1260 11462
rect 980 10332 1036 10342
rect 980 10108 1036 10276
rect 1204 10332 1260 11396
rect 1204 10266 1260 10276
rect 1316 11228 1372 11238
rect 980 10042 1036 10052
rect 868 9818 924 9828
rect 1092 9884 1148 9894
rect 644 9772 700 9782
rect 644 9553 700 9716
rect 980 9772 1036 9782
rect 756 9553 812 9563
rect 644 9497 756 9553
rect 756 9487 812 9497
rect 644 9426 700 9436
rect 700 9370 812 9426
rect 644 9360 700 9370
rect 308 8586 364 8596
rect 756 9299 812 9309
rect 84 8428 140 8438
rect 140 8372 252 8428
rect 84 8362 140 8372
rect 84 4956 140 5068
rect 84 4890 140 4900
rect 84 4732 140 4742
rect 84 4172 140 4676
rect 84 4106 140 4116
rect 196 1372 252 8372
rect 420 5180 476 5190
rect 420 4956 476 5124
rect 420 4890 476 4900
rect 308 4396 364 4406
rect 308 4284 364 4340
rect 756 4396 812 9243
rect 980 9304 1036 9716
rect 980 9238 1036 9248
rect 980 8764 1036 8774
rect 980 8652 1036 8708
rect 980 8586 1036 8596
rect 1092 8540 1148 9828
rect 1316 9772 1372 11172
rect 1316 9706 1372 9716
rect 1428 10332 1484 13860
rect 1540 13244 1596 14308
rect 1652 14140 1708 14868
rect 1876 14364 1932 16548
rect 2212 16589 2268 16660
rect 2324 16716 2380 16828
rect 2324 16650 2380 16660
rect 2436 16716 2492 16884
rect 2548 16828 2604 17444
rect 2660 17714 2716 17724
rect 2660 17500 2716 17658
rect 2660 17434 2716 17444
rect 2548 16772 2558 16828
rect 2614 16772 2624 16828
rect 2884 16716 2940 16726
rect 2436 16650 2492 16660
rect 2548 16701 2604 16711
rect 2548 16533 2604 16645
rect 2884 16609 2940 16660
rect 2884 16543 2940 16553
rect 2212 16523 2268 16533
rect 2772 16492 2828 16502
rect 2772 15820 2828 16436
rect 2772 15754 2828 15764
rect 2884 16472 2940 16482
rect 2884 15820 2940 16416
rect 2548 15708 2604 15718
rect 1988 15148 2044 15158
rect 1988 14980 2044 15092
rect 2436 15036 2492 15046
rect 2436 14924 2492 14980
rect 2436 14858 2492 14868
rect 1876 14298 1932 14308
rect 2548 14700 2604 15652
rect 2884 15596 2940 15764
rect 2996 15708 3052 19348
rect 3332 20300 3388 20356
rect 4004 20320 4060 20330
rect 4116 20320 4172 20468
rect 3108 18396 3164 18406
rect 3108 18080 3164 18340
rect 3332 18396 3388 20244
rect 3668 20300 3724 20310
rect 3668 20076 3724 20244
rect 3780 20188 3836 20300
rect 4060 20264 4172 20320
rect 4340 20300 4396 20310
rect 4004 20254 4060 20264
rect 3780 20122 3836 20132
rect 4116 20188 4172 20198
rect 4172 20132 4284 20188
rect 4116 20122 4172 20132
rect 3668 20010 3724 20020
rect 4228 20056 4284 20066
rect 4228 19628 4284 20000
rect 4228 19562 4284 19572
rect 3892 19292 3948 19302
rect 3892 19180 3948 19236
rect 3444 19068 3500 19078
rect 3444 18508 3500 19012
rect 3444 18442 3500 18452
rect 3668 18508 3724 18518
rect 3332 18330 3388 18340
rect 3668 18396 3724 18452
rect 3668 18330 3724 18340
rect 3780 18508 3836 18518
rect 3240 18172 3296 18182
rect 3108 18014 3164 18024
rect 3220 18116 3240 18172
rect 3220 18106 3296 18116
rect 3780 18172 3836 18452
rect 3780 18106 3836 18116
rect 3892 18508 3948 19124
rect 4116 19292 4172 19302
rect 4116 18732 4172 19236
rect 4116 18666 4172 18676
rect 3108 17943 3164 17953
rect 3108 17500 3164 17887
rect 3108 17434 3164 17444
rect 3220 17500 3276 18106
rect 3220 17434 3276 17444
rect 3556 17500 3612 17612
rect 3556 17434 3612 17444
rect 3668 17500 3724 17510
rect 3108 17276 3164 17286
rect 3108 16726 3164 17220
rect 3230 17276 3286 17286
rect 3230 17164 3286 17220
rect 3230 17098 3286 17108
rect 3525 16772 3536 16828
rect 3592 16772 3612 16828
rect 3108 16660 3164 16670
rect 3556 16716 3612 16772
rect 3556 16650 3612 16660
rect 3668 16716 3724 17444
rect 3892 17276 3948 18452
rect 4116 18284 4172 18294
rect 4116 17948 4172 18228
rect 4116 17882 4172 17892
rect 4228 17612 4284 17622
rect 4116 17500 4172 17612
rect 4228 17444 4284 17556
rect 4116 17434 4172 17444
rect 3892 17119 3948 17220
rect 3534 16538 3544 16594
rect 3600 16538 3610 16594
rect 3544 16482 3600 16538
rect 3544 16428 3612 16482
rect 3556 16380 3612 16428
rect 3556 16314 3612 16324
rect 3108 15820 3164 15932
rect 3108 15754 3164 15764
rect 2996 15642 3052 15652
rect 2884 15530 2940 15540
rect 3220 15148 3276 15158
rect 1652 14074 1708 14084
rect 2548 13916 2604 14644
rect 2660 14924 2716 14934
rect 2660 14476 2716 14868
rect 3220 14924 3276 15092
rect 3668 15036 3724 16660
rect 3668 14970 3724 14980
rect 3780 17063 3948 17119
rect 3780 16716 3836 17063
rect 4340 17052 4396 20244
rect 4452 20300 4508 20412
rect 4452 20234 4508 20244
rect 4676 20300 4732 20310
rect 5012 20300 5068 20310
rect 4900 20244 5012 20300
rect 4676 20188 4732 20244
rect 5012 20234 5068 20244
rect 5348 20300 5404 20310
rect 6020 20300 6076 20310
rect 5908 20244 6020 20300
rect 5348 20132 5404 20244
rect 6020 20234 6076 20244
rect 6356 20300 6412 20310
rect 6356 20132 6412 20244
rect 7364 20300 7420 20310
rect 4452 19516 4508 19526
rect 4452 19292 4508 19460
rect 4452 19226 4508 19236
rect 4564 19292 4620 19302
rect 4564 19180 4620 19236
rect 4564 19114 4620 19124
rect 4340 16986 4396 16996
rect 4452 18956 4508 18966
rect 4452 18508 4508 18900
rect 4676 18844 4732 20132
rect 4900 20076 4956 20086
rect 4900 19516 4956 20020
rect 6244 20076 6300 20086
rect 6244 19964 6300 20020
rect 6244 19898 6300 19908
rect 5992 19740 6044 19796
rect 6100 19740 6200 19796
rect 6256 19740 6356 19796
rect 6412 19740 6512 19796
rect 6568 19740 6668 19796
rect 6724 19740 6776 19796
rect 4900 19450 4956 19460
rect 4788 19312 4844 19322
rect 4844 19256 4956 19312
rect 5348 19292 5404 19302
rect 4788 19246 4844 19256
rect 4788 19180 4844 19190
rect 4788 19068 4844 19124
rect 4788 19002 4844 19012
rect 5124 19180 5180 19190
rect 4676 18778 4732 18788
rect 4900 18844 4956 18854
rect 4900 18732 4956 18788
rect 4900 18666 4956 18676
rect 3220 14858 3276 14868
rect 3780 14924 3836 16660
rect 3892 16828 3948 16838
rect 3892 16716 3948 16772
rect 4228 16828 4284 16838
rect 4116 16716 4172 16726
rect 4004 16660 4116 16716
rect 4228 16660 4284 16772
rect 4452 16716 4508 18452
rect 4676 18508 4732 18518
rect 4676 18396 4732 18452
rect 5124 18508 5180 19124
rect 5348 19068 5404 19236
rect 5348 19002 5404 19012
rect 7140 19180 7196 19190
rect 7140 19068 7196 19124
rect 7140 19002 7196 19012
rect 6468 18956 6524 18966
rect 5796 18620 5852 18732
rect 5796 18554 5852 18564
rect 4676 18330 4732 18340
rect 4900 18396 4956 18406
rect 4564 18284 4620 18294
rect 4564 18172 4620 18228
rect 4900 18284 4956 18340
rect 4900 18218 4956 18228
rect 4564 18106 4620 18116
rect 5124 17500 5180 18452
rect 5236 18508 5292 18518
rect 5236 18284 5292 18452
rect 5236 17724 5292 18228
rect 5572 18508 5628 18518
rect 5572 18284 5628 18452
rect 5572 18218 5628 18228
rect 5684 18508 5740 18518
rect 5236 17658 5292 17668
rect 5124 17434 5180 17444
rect 5684 17052 5740 18452
rect 6132 18508 6188 18518
rect 5908 18396 5964 18406
rect 5796 18340 5908 18396
rect 5908 18330 5964 18340
rect 6132 18284 6188 18452
rect 6244 18508 6300 18620
rect 6244 18441 6300 18452
rect 6356 18508 6412 18620
rect 6356 18442 6412 18452
rect 6468 18508 6524 18900
rect 7364 18732 7420 20244
rect 8820 20300 8876 20310
rect 8820 20188 8876 20244
rect 10276 20300 10332 20310
rect 8820 20122 8876 20132
rect 9044 20188 9100 20198
rect 7364 18666 7420 18676
rect 8036 19292 8092 19302
rect 6468 18442 6524 18452
rect 7588 18620 7644 18630
rect 7588 18508 7644 18564
rect 7588 18442 7644 18452
rect 7700 18508 7756 18518
rect 6132 18218 6188 18228
rect 7364 18396 7420 18406
rect 7700 18340 7756 18452
rect 8036 18508 8092 19236
rect 9044 19292 9100 20132
rect 9380 19964 9436 19974
rect 9044 19226 9100 19236
rect 9156 19404 9212 19414
rect 5992 17948 6044 18004
rect 6100 17948 6200 18004
rect 6256 17948 6356 18004
rect 6412 17948 6512 18004
rect 6568 17948 6668 18004
rect 6724 17948 6776 18004
rect 5684 16986 5740 16996
rect 6804 17612 6860 17622
rect 5460 16940 5516 16950
rect 3892 16650 3948 16660
rect 4116 16650 4172 16660
rect 4452 16650 4508 16660
rect 4564 16716 4620 16726
rect 5460 16716 5516 16884
rect 4564 16604 4620 16660
rect 4564 16538 4620 16548
rect 5348 16604 5404 16716
rect 5348 16538 5404 16548
rect 4340 15932 4396 15942
rect 4228 15596 4284 15606
rect 3780 14858 3836 14868
rect 4004 15036 4060 15046
rect 2660 14410 2716 14420
rect 2772 14812 2828 14822
rect 2548 13850 2604 13860
rect 1876 13804 1932 13814
rect 1876 13356 1932 13748
rect 1876 13290 1932 13300
rect 2324 13468 2380 13478
rect 1540 13178 1596 13188
rect 2212 13132 2268 13142
rect 1764 13020 1820 13030
rect 1820 12964 1932 13020
rect 1764 12954 1820 12964
rect 1876 12348 1932 12358
rect 1652 11228 1708 11238
rect 1652 11060 1708 11172
rect 1876 11228 1932 12292
rect 2212 12124 2268 13076
rect 2324 13132 2380 13412
rect 2324 13066 2380 13076
rect 2772 13356 2828 14756
rect 3108 14812 3164 14822
rect 3108 14145 3164 14756
rect 3780 14700 3836 14710
rect 3836 14644 3948 14700
rect 3780 14634 3836 14644
rect 3892 14252 3948 14644
rect 3108 14079 3164 14089
rect 3332 14140 3388 14150
rect 3332 14028 3388 14084
rect 3108 13916 3164 14015
rect 3332 13962 3388 13972
rect 3892 14028 3948 14196
rect 3892 13962 3948 13972
rect 3108 13850 3164 13860
rect 3668 13916 3724 13926
rect 2996 13804 3052 13814
rect 2996 13468 3052 13748
rect 2996 13402 3052 13412
rect 2436 13020 2492 13030
rect 2492 12964 2604 13020
rect 2436 12954 2492 12964
rect 2212 12058 2268 12068
rect 2436 12124 2492 12134
rect 2436 11340 2492 12068
rect 2436 11274 2492 11284
rect 1428 9660 1484 10276
rect 1652 10332 1708 10342
rect 1708 10276 1820 10332
rect 1652 10266 1708 10276
rect 1876 10220 1932 11172
rect 2324 10332 2380 10342
rect 2380 10276 2492 10332
rect 2324 10266 2380 10276
rect 1876 10154 1932 10164
rect 1652 10108 1708 10118
rect 1428 9594 1484 9604
rect 1204 9548 1260 9558
rect 1540 9538 1596 9660
rect 1204 8876 1260 9492
rect 1510 9482 1520 9538
rect 1652 9558 1708 10052
rect 2548 9772 2604 12964
rect 2772 10664 2828 13300
rect 3444 13356 3500 13366
rect 3332 13132 3388 13244
rect 2996 12796 3052 12806
rect 2884 12740 2996 12796
rect 2996 12730 3052 12740
rect 3220 12124 3276 12236
rect 3220 12058 3276 12068
rect 2996 11340 3052 11350
rect 2996 10892 3052 11284
rect 2996 10826 3052 10836
rect 3332 10668 3388 13076
rect 3444 13132 3500 13300
rect 3668 13356 3724 13860
rect 3668 13290 3724 13300
rect 4004 13916 4060 14980
rect 4116 14924 4172 14934
rect 4228 14924 4284 15540
rect 4172 14868 4284 14924
rect 4116 14858 4172 14868
rect 4228 14140 4284 14868
rect 4228 14028 4284 14084
rect 4340 14140 4396 15876
rect 4564 15708 4620 15718
rect 4564 15596 4620 15652
rect 4564 15061 4620 15540
rect 4900 15708 4956 15718
rect 4900 15596 4956 15652
rect 4788 15260 4844 15270
rect 4788 15148 4844 15204
rect 4788 15082 4844 15092
rect 4452 15051 4620 15061
rect 4508 14995 4620 15051
rect 4452 14985 4508 14995
rect 4564 14924 4620 14934
rect 4452 14868 4564 14924
rect 4620 14868 4732 14924
rect 4564 14858 4620 14868
rect 4340 14074 4396 14084
rect 4564 14476 4620 14486
rect 4218 13972 4228 14028
rect 4284 13972 4294 14028
rect 4564 13916 4620 14420
rect 3444 13066 3500 13076
rect 4004 13132 4060 13860
rect 4228 13906 4284 13916
rect 4004 13066 4060 13076
rect 4116 13356 4172 13366
rect 4116 13132 4172 13300
rect 3556 12236 3612 12246
rect 3612 12180 3724 12236
rect 3556 12170 3612 12180
rect 3892 12124 3948 12236
rect 3892 12058 3948 12068
rect 4116 12124 4172 13076
rect 4228 13356 4284 13850
rect 4228 12460 4284 13300
rect 4340 13692 4396 13702
rect 4340 13132 4396 13636
rect 4564 13356 4620 13860
rect 4676 13916 4732 14868
rect 4676 13692 4732 13860
rect 4788 14812 4844 14822
rect 4788 13916 4844 14756
rect 4900 14476 4956 15540
rect 5348 15708 5404 15718
rect 5348 15596 5404 15652
rect 5348 15530 5404 15540
rect 4900 14410 4956 14420
rect 5236 15372 5292 15382
rect 4900 14252 4956 14262
rect 4900 14028 4956 14196
rect 4900 13962 4956 13972
rect 5236 14028 5292 15316
rect 5460 15372 5516 16660
rect 5908 16716 5964 16828
rect 5908 16650 5964 16660
rect 6020 16716 6076 16726
rect 5796 16604 5852 16614
rect 5684 16548 5796 16604
rect 5796 16538 5852 16548
rect 5796 16380 5852 16390
rect 5796 16044 5852 16324
rect 6020 16380 6076 16660
rect 6804 16492 6860 17556
rect 6804 16426 6860 16436
rect 7028 17612 7084 17622
rect 7028 16492 7084 17556
rect 7364 17612 7420 18340
rect 7364 17546 7420 17556
rect 7588 16828 7644 16838
rect 7364 16716 7420 16726
rect 7252 16660 7364 16716
rect 7364 16650 7420 16660
rect 7588 16716 7644 16772
rect 7588 16650 7644 16660
rect 7700 16716 7756 16726
rect 7242 16543 7252 16599
rect 7308 16543 7318 16599
rect 7028 16426 7084 16436
rect 6020 16314 6076 16324
rect 5992 16156 6044 16212
rect 6100 16156 6200 16212
rect 6256 16156 6356 16212
rect 6412 16156 6512 16212
rect 6568 16156 6668 16212
rect 6724 16156 6776 16212
rect 5796 15978 5852 15988
rect 6356 16044 6412 16054
rect 6356 15927 6412 15988
rect 6346 15871 6356 15927
rect 6412 15871 6422 15927
rect 7252 15820 7308 16543
rect 5572 15708 5628 15820
rect 5572 15642 5628 15652
rect 5796 15708 5852 15718
rect 5460 15306 5516 15316
rect 5796 15372 5852 15652
rect 6020 15708 6076 15718
rect 6020 15596 6076 15652
rect 6132 15708 6188 15820
rect 6132 15642 6188 15652
rect 6356 15805 6412 15815
rect 7252 15754 7308 15764
rect 7588 15932 7644 15942
rect 7700 15932 7756 16660
rect 7644 15876 7756 15932
rect 7812 16716 7868 16726
rect 7812 15932 7868 16660
rect 6356 15708 6412 15749
rect 7364 15708 7420 15718
rect 6020 15530 6076 15540
rect 5796 14252 5852 15316
rect 6356 14924 6412 15652
rect 6468 15688 6524 15698
rect 6468 15036 6524 15632
rect 7364 15382 7420 15652
rect 7588 15708 7644 15876
rect 7812 15866 7868 15876
rect 7924 16716 7980 16726
rect 7588 15642 7644 15652
rect 7344 15372 7420 15382
rect 7481 15372 7537 15382
rect 7400 15316 7420 15372
rect 7476 15316 7481 15372
rect 7344 15306 7400 15316
rect 7476 15306 7537 15316
rect 7924 15372 7980 16660
rect 7924 15306 7980 15316
rect 6468 14970 6524 14980
rect 6356 14858 6412 14868
rect 7252 14924 7308 14934
rect 6804 14700 6860 14710
rect 6804 14588 6860 14644
rect 7252 14700 7308 14868
rect 7252 14634 7308 14644
rect 6804 14522 6860 14532
rect 5992 14364 6044 14420
rect 6100 14364 6200 14420
rect 6256 14364 6356 14420
rect 6412 14364 6512 14420
rect 6568 14364 6668 14420
rect 6724 14364 6776 14420
rect 5796 14186 5852 14196
rect 6132 14252 6188 14262
rect 6132 14140 6188 14196
rect 6132 14074 6188 14084
rect 7476 14140 7532 15306
rect 8036 14700 8092 18452
rect 8148 18396 8204 18406
rect 8932 18396 8988 18406
rect 8148 16716 8204 18340
rect 8820 18340 8932 18396
rect 8148 15484 8204 16660
rect 8260 17500 8316 17510
rect 8260 15708 8316 17444
rect 8820 16940 8876 18340
rect 8932 18330 8988 18340
rect 9156 18396 9212 19348
rect 9380 19404 9436 19908
rect 9380 19338 9436 19348
rect 10276 19180 10332 20244
rect 11956 20300 12012 20412
rect 11956 20234 12012 20244
rect 12292 20300 12348 20310
rect 10948 20188 11004 20198
rect 11004 20132 11116 20188
rect 10948 20122 11004 20132
rect 12292 19852 12348 20244
rect 12740 20188 12796 20198
rect 12740 20020 12796 20132
rect 13076 20188 13132 20972
rect 16408 20636 16460 20692
rect 16516 20636 16616 20692
rect 16672 20636 16772 20692
rect 16828 20636 16928 20692
rect 16984 20636 17084 20692
rect 17140 20636 17192 20692
rect 20468 20412 20524 20422
rect 14084 20300 14140 20310
rect 12292 19786 12348 19796
rect 12852 19964 12908 19974
rect 10276 19114 10332 19124
rect 10388 19404 10444 19414
rect 10276 18508 10332 18518
rect 10164 18452 10276 18508
rect 10276 18442 10332 18452
rect 8820 16874 8876 16884
rect 9044 17388 9100 17500
rect 9044 16828 9100 17332
rect 8372 16716 8433 16726
rect 8372 16650 8433 16660
rect 8489 16716 8565 16726
rect 8932 16716 8988 16828
rect 8565 16660 8652 16716
rect 8489 16650 8565 16660
rect 8932 16650 8988 16660
rect 9044 16716 9100 16772
rect 9044 16650 9100 16660
rect 8377 16604 8433 16650
rect 8377 16538 8433 16548
rect 8260 15642 8316 15652
rect 8484 16492 8540 16502
rect 8148 15418 8204 15428
rect 8036 14634 8092 14644
rect 8372 14812 8428 14822
rect 4788 13850 4844 13860
rect 4676 13626 4732 13636
rect 4564 13290 4620 13300
rect 4340 13066 4396 13076
rect 4452 13244 4508 13254
rect 4228 12394 4284 12404
rect 4340 12796 4396 12806
rect 4004 11340 4060 11350
rect 2752 10595 2828 10664
rect 3220 10612 3388 10668
rect 3780 11228 3836 11238
rect 2752 10444 2808 10595
rect 2752 10378 2808 10388
rect 2864 10444 2920 10454
rect 2996 10444 3057 10454
rect 2920 10388 2940 10444
rect 2864 10378 2940 10388
rect 3057 10388 3164 10444
rect 2996 10378 3057 10388
rect 2548 9706 2604 9716
rect 1652 9548 1713 9558
rect 1871 9548 1932 9558
rect 1652 9492 1657 9548
rect 1780 9492 1871 9548
rect 1657 9482 1713 9492
rect 1871 9482 1932 9492
rect 1988 9548 2064 9558
rect 2212 9548 2268 9558
rect 2064 9492 2156 9548
rect 1988 9482 2064 9492
rect 1540 9472 1596 9482
rect 1204 8810 1260 8820
rect 756 4330 812 4340
rect 868 6860 924 6870
rect 868 4396 924 6804
rect 1092 5292 1148 8484
rect 1876 7644 1932 7756
rect 1876 7578 1932 7588
rect 2100 7644 2156 7654
rect 1876 6860 1932 6870
rect 2100 6860 2156 7588
rect 1876 6692 1932 6804
rect 1988 6804 2100 6860
rect 1652 6076 1708 6086
rect 1652 5852 1708 6020
rect 1652 5786 1708 5796
rect 1876 5852 1932 5862
rect 1988 5852 2044 6804
rect 2100 6794 2156 6804
rect 1932 5796 2044 5852
rect 1876 5786 1932 5796
rect 1092 5226 1148 5236
rect 1428 5292 1484 5302
rect 1092 4956 1148 5068
rect 1092 4890 1148 4900
rect 868 4330 924 4340
rect 1316 4508 1372 4518
rect 308 4218 364 4228
rect 420 4172 476 4182
rect 980 4172 1036 4284
rect 476 4116 588 4172
rect 420 4106 476 4116
rect 980 4106 1036 4116
rect 1316 4172 1372 4452
rect 868 3276 924 3388
rect 868 3210 924 3220
rect 1316 3276 1372 4116
rect 1316 3210 1372 3220
rect 1428 3388 1484 5236
rect 1540 5068 1596 5078
rect 1540 4956 1596 5012
rect 1540 4890 1596 4900
rect 1764 4956 1820 4966
rect 1764 4732 1820 4900
rect 1876 4956 1932 5068
rect 1876 4890 1932 4900
rect 1764 4666 1820 4676
rect 1988 4712 2044 5796
rect 2100 4956 2156 4966
rect 2100 4844 2156 4900
rect 2100 4778 2156 4788
rect 2212 4956 2268 9492
rect 2548 9487 2660 9543
rect 2716 9487 2726 9543
rect 2324 9324 2380 9334
rect 2324 8652 2380 9268
rect 2548 8764 2604 9487
rect 2660 9421 2716 9431
rect 2716 9365 2828 9421
rect 2660 9355 2716 9365
rect 2548 8698 2604 8708
rect 2884 8764 2940 10378
rect 3220 10332 3276 10612
rect 3220 10266 3276 10276
rect 3332 10332 3388 10444
rect 3332 10266 3388 10276
rect 3556 10220 3612 10230
rect 3332 10108 3388 10118
rect 3220 9284 3276 9294
rect 2884 8698 2940 8708
rect 2324 8586 2380 8596
rect 2436 8652 2492 8662
rect 2436 8540 2492 8596
rect 2996 8652 3052 8764
rect 2996 8586 3052 8596
rect 2324 5180 2380 5190
rect 2324 5012 2380 5124
rect 2436 5068 2492 8484
rect 2660 8540 2716 8550
rect 2660 7873 2716 8484
rect 2660 7807 2716 7817
rect 2772 8540 2828 8550
rect 2212 4732 2268 4900
rect 2436 4956 2492 5012
rect 2436 4890 2492 4900
rect 2660 7736 2716 7746
rect 2660 4956 2716 7680
rect 2772 5068 2828 8484
rect 3108 8540 3164 8550
rect 3220 8540 3276 9228
rect 3164 8484 3276 8540
rect 3332 8540 3388 10052
rect 3444 9548 3500 9558
rect 3444 9436 3500 9492
rect 3444 9370 3500 9380
rect 3556 8896 3612 10164
rect 3668 10220 3724 10230
rect 3668 9884 3724 10164
rect 3668 9818 3724 9828
rect 3780 9548 3836 11172
rect 3780 9482 3836 9492
rect 3892 9772 3948 9782
rect 3892 9553 3948 9716
rect 3892 9487 3948 9497
rect 3556 8830 3612 8840
rect 3668 9436 3724 9446
rect 3556 8759 3612 8769
rect 3556 8652 3612 8703
rect 3556 8586 3612 8596
rect 3108 8474 3164 8484
rect 3332 8474 3388 8484
rect 3444 8428 3500 8438
rect 3444 8092 3500 8372
rect 3444 8026 3500 8036
rect 3556 8316 3612 8326
rect 3444 7868 3500 7878
rect 3220 7756 3276 7766
rect 3220 6748 3276 7700
rect 3108 6692 3220 6748
rect 2772 5002 2828 5012
rect 2884 6188 2940 6198
rect 2884 5068 2940 6132
rect 3108 5964 3164 6692
rect 3220 6682 3276 6692
rect 2660 4890 2716 4900
rect 2884 4844 2940 5012
rect 2996 5068 3052 5078
rect 2996 4956 3052 5012
rect 2996 4890 3052 4900
rect 2884 4778 2940 4788
rect 3108 4824 3164 5908
rect 3332 5292 3388 5302
rect 3220 5068 3276 5078
rect 3220 4956 3276 5012
rect 3220 4890 3276 4900
rect 3332 4956 3388 5236
rect 3332 4890 3388 4900
rect 3444 5180 3500 7812
rect 3556 7644 3612 8260
rect 3556 7578 3612 7588
rect 3668 7512 3724 9380
rect 3780 9411 3836 9421
rect 3836 9355 3948 9411
rect 3780 9345 3836 9355
rect 3780 8876 3836 8886
rect 3780 8540 3836 8820
rect 3780 8474 3836 8484
rect 3892 8540 3948 8550
rect 3892 8316 3948 8484
rect 3892 8250 3948 8260
rect 4004 8428 4060 11284
rect 4116 11228 4172 12068
rect 4340 11340 4396 12740
rect 4340 11274 4396 11284
rect 4452 12236 4508 13188
rect 5236 13244 5292 13972
rect 5572 14028 5628 14038
rect 5236 13178 5292 13188
rect 5460 13692 5516 13702
rect 4676 13132 4732 13142
rect 4564 12908 4620 12918
rect 4564 12460 4620 12852
rect 4564 12394 4620 12404
rect 4676 12348 4732 13076
rect 4676 12282 4732 12292
rect 5348 12348 5404 12358
rect 4116 10444 4172 11172
rect 4116 10378 4172 10388
rect 4452 10108 4508 12180
rect 5236 12012 5292 12022
rect 5236 11452 5292 11956
rect 5348 12012 5404 12292
rect 5348 11946 5404 11956
rect 5236 11386 5292 11396
rect 4676 11340 4732 11350
rect 4564 11228 4620 11340
rect 4732 11284 4844 11340
rect 4676 11274 4732 11284
rect 4564 11162 4620 11172
rect 4778 11167 4788 11223
rect 4844 11167 4854 11223
rect 4788 10892 4844 11167
rect 4788 10332 4844 10836
rect 5236 11116 5292 11126
rect 5236 10444 5292 11060
rect 5236 10378 5292 10388
rect 4788 10266 4844 10276
rect 4452 10042 4508 10052
rect 4116 9660 4172 9670
rect 4116 9548 4172 9604
rect 4452 9660 4508 9670
rect 4116 9482 4172 9492
rect 4228 9416 4284 9548
rect 4228 9350 4284 9360
rect 4116 8876 4172 8886
rect 4116 8550 4172 8820
rect 4116 8484 4172 8494
rect 4452 8540 4508 9604
rect 4676 9548 4732 9558
rect 4676 9324 4732 9492
rect 4676 9258 4732 9268
rect 4340 8483 4396 8493
rect 3444 4956 3500 5124
rect 3444 4890 3500 4900
rect 3556 7456 3724 7512
rect 3892 8092 3948 8102
rect 3108 4768 3276 4824
rect 1988 4656 2156 4712
rect 2212 4666 2268 4676
rect 2548 4732 2604 4742
rect 1876 4620 1932 4630
rect 1540 4284 1596 4294
rect 1540 4172 1596 4228
rect 1540 4106 1596 4116
rect 1652 4172 1708 4182
rect 1876 4172 1932 4564
rect 1708 4116 1820 4172
rect 1652 4106 1708 4116
rect 308 3052 364 3062
rect 308 1484 364 2996
rect 644 3052 700 3062
rect 644 2884 700 2996
rect 1428 1596 1484 3332
rect 1540 3276 1596 3388
rect 1540 3210 1596 3220
rect 1876 3276 1932 4116
rect 1988 4172 2044 4182
rect 1988 3948 2044 4116
rect 1988 3882 2044 3892
rect 1876 3210 1932 3220
rect 1876 2940 1932 2950
rect 1652 2716 1708 2726
rect 1876 2721 1932 2884
rect 1866 2665 1876 2721
rect 1932 2665 1942 2721
rect 1652 2268 1708 2660
rect 1652 2202 1708 2212
rect 1876 2599 1932 2609
rect 1876 2268 1932 2543
rect 2100 2604 2156 4656
rect 2436 4284 2492 4294
rect 2324 4172 2380 4284
rect 2212 4060 2268 4172
rect 2324 4106 2380 4116
rect 2212 3994 2268 4004
rect 2212 3276 2268 3286
rect 2268 3220 2380 3276
rect 2212 3210 2268 3220
rect 2436 3164 2492 4228
rect 2548 3388 2604 4676
rect 2884 4396 2940 4508
rect 2884 4330 2940 4340
rect 2772 4284 2828 4294
rect 2660 4172 2716 4182
rect 2660 4060 2716 4116
rect 2660 3994 2716 4004
rect 2548 3322 2604 3332
rect 2436 3098 2492 3108
rect 2548 3164 2604 3174
rect 2772 3164 2828 4228
rect 3108 4172 3164 4182
rect 3108 4060 3164 4116
rect 3108 3994 3164 4004
rect 3220 3928 3276 4768
rect 3108 3872 3276 3928
rect 2604 3108 2716 3164
rect 2548 3098 2604 3108
rect 2772 3098 2828 3108
rect 2996 3164 3052 3174
rect 2100 2538 2156 2548
rect 1428 1530 1484 1540
rect 1764 1708 1820 1718
rect 308 1418 364 1428
rect 868 1484 924 1494
rect 196 1306 252 1316
rect 868 812 924 1428
rect 1204 1484 1260 1494
rect 1204 1372 1260 1428
rect 1764 1484 1820 1652
rect 1764 1418 1820 1428
rect 1204 1306 1260 1316
rect 868 746 924 756
rect 1652 1036 1708 1046
rect 1652 476 1708 980
rect 1652 410 1708 420
rect 1876 476 1932 2212
rect 2324 1596 2380 1708
rect 2324 1530 2380 1540
rect 2436 1484 2492 1494
rect 2996 1484 3052 3108
rect 2492 1428 2604 1484
rect 2436 1418 2492 1428
rect 2996 1418 3052 1428
rect 3108 2380 3164 3872
rect 3444 3276 3500 3388
rect 3444 3210 3500 3220
rect 3556 2828 3612 7456
rect 3892 6860 3948 8036
rect 4004 7756 4060 8372
rect 4116 8316 4172 8428
rect 4228 8372 4340 8428
rect 4340 8362 4396 8372
rect 4116 8250 4172 8260
rect 4004 7690 4060 7700
rect 4452 7756 4508 8484
rect 5460 8652 5516 13636
rect 5572 12460 5628 13972
rect 6244 14028 6300 14038
rect 5796 13916 5852 13926
rect 5796 13249 5852 13860
rect 6244 13916 6300 13972
rect 6244 13850 6300 13860
rect 7364 13916 7420 13926
rect 7364 13748 7420 13860
rect 7476 13916 7532 14084
rect 7924 14588 7980 14598
rect 7924 14028 7980 14532
rect 7924 13962 7980 13972
rect 8148 14140 8204 14150
rect 7476 13850 7532 13860
rect 7700 13916 7756 13926
rect 5796 13183 5852 13193
rect 6020 13692 6076 13702
rect 5786 13071 5796 13127
rect 5852 13071 5862 13127
rect 5572 12394 5628 12404
rect 5684 12124 5740 12134
rect 5572 12068 5684 12124
rect 5684 12058 5740 12068
rect 5796 12124 5852 13071
rect 6020 13020 6076 13636
rect 7700 13692 7756 13860
rect 7700 13626 7756 13636
rect 7812 13916 7868 13926
rect 6020 12954 6076 12964
rect 7140 13020 7196 13132
rect 7364 13020 7420 13030
rect 7140 12954 7196 12964
rect 7252 12964 7364 13020
rect 5992 12572 6044 12628
rect 6100 12572 6200 12628
rect 6256 12572 6356 12628
rect 6412 12572 6512 12628
rect 6568 12572 6668 12628
rect 6724 12572 6776 12628
rect 5796 12058 5852 12068
rect 6916 12348 6972 12358
rect 6916 12124 6972 12292
rect 6244 11900 6300 11910
rect 6244 11788 6300 11844
rect 6244 11722 6300 11732
rect 6916 11228 6972 12068
rect 6916 11162 6972 11172
rect 5992 10780 6044 10836
rect 6100 10780 6200 10836
rect 6256 10780 6356 10836
rect 6412 10780 6512 10836
rect 6568 10780 6668 10836
rect 6724 10780 6776 10836
rect 6020 10444 6076 10454
rect 6020 10220 6076 10388
rect 6244 10444 6300 10556
rect 6244 10378 6300 10388
rect 6020 10154 6076 10164
rect 6804 10220 6860 10230
rect 5684 9436 5740 9446
rect 5684 8764 5740 9380
rect 6580 9436 6636 9446
rect 6580 9268 6636 9380
rect 6804 9436 6860 10164
rect 7252 10220 7308 12964
rect 7364 12954 7420 12964
rect 7588 12246 7644 12256
rect 7476 12124 7532 12134
rect 7364 12068 7476 12124
rect 7588 12068 7644 12190
rect 7812 12134 7868 13860
rect 8036 12460 8092 12470
rect 8036 12236 8092 12404
rect 8036 12170 8092 12180
rect 7868 12078 7980 12134
rect 7812 12068 7868 12078
rect 7476 12058 7532 12068
rect 7700 12012 7756 12022
rect 7756 11956 7868 12012
rect 7924 12007 7980 12017
rect 7700 11946 7756 11956
rect 7924 11844 7980 11951
rect 7700 11340 7756 11350
rect 7700 11228 7756 11284
rect 7700 11162 7756 11172
rect 7924 11228 7980 11238
rect 7252 10154 7308 10164
rect 7924 9548 7980 11172
rect 7924 9482 7980 9492
rect 6804 9370 6860 9380
rect 5992 8988 6044 9044
rect 6100 8988 6200 9044
rect 6256 8988 6356 9044
rect 6412 8988 6512 9044
rect 6568 8988 6668 9044
rect 6724 8988 6776 9044
rect 8148 8876 8204 14084
rect 8372 14140 8428 14756
rect 8484 14812 8540 16436
rect 9156 16492 9212 18340
rect 9380 17500 9436 17510
rect 9716 17500 9772 17510
rect 9436 17444 9548 17500
rect 9380 17388 9436 17444
rect 9380 17322 9436 17332
rect 9492 16940 9548 17444
rect 9716 17388 9772 17444
rect 9716 17322 9772 17332
rect 9940 17388 9996 17398
rect 9940 17276 9996 17332
rect 9940 17210 9996 17220
rect 9268 16716 9324 16726
rect 9268 16604 9324 16660
rect 9492 16609 9548 16884
rect 9716 16726 9772 16736
rect 9940 16726 9996 16736
rect 9772 16670 9884 16726
rect 9716 16660 9772 16670
rect 9482 16553 9492 16609
rect 9548 16553 9558 16609
rect 9828 16599 9884 16609
rect 9268 16538 9324 16548
rect 9156 16426 9212 16436
rect 9492 16487 9548 16497
rect 9268 15820 9324 15932
rect 9268 15754 9324 15764
rect 9492 15820 9548 16431
rect 9492 15754 9548 15764
rect 9716 16492 9772 16502
rect 8708 14812 8764 14822
rect 8596 14756 8708 14812
rect 8484 14746 8540 14756
rect 8708 14746 8764 14756
rect 9380 14252 9436 14262
rect 9268 14196 9380 14252
rect 9380 14186 9436 14196
rect 8372 14074 8428 14084
rect 9044 13916 9100 13926
rect 8820 13804 8876 13814
rect 8372 13692 8428 13702
rect 8372 12236 8428 13636
rect 8372 12170 8428 12180
rect 8484 13132 8540 13142
rect 8484 11228 8540 13076
rect 8820 12796 8876 13748
rect 9044 13244 9100 13860
rect 9492 13916 9548 13926
rect 9380 13692 9436 13804
rect 9380 13626 9436 13636
rect 9044 13178 9100 13188
rect 8708 12348 8764 12358
rect 8596 12236 8652 12246
rect 8596 12124 8652 12180
rect 8596 12058 8652 12068
rect 8484 11162 8540 11172
rect 8708 11228 8764 12292
rect 8820 12348 8876 12740
rect 8820 12282 8876 12292
rect 9268 12908 9324 12918
rect 9268 12572 9324 12852
rect 9044 12124 9100 12134
rect 9044 11340 9100 12068
rect 9156 12124 9212 12236
rect 9156 12058 9212 12068
rect 8708 11162 8764 11172
rect 8932 11228 8988 11238
rect 8932 10220 8988 11172
rect 8932 10154 8988 10164
rect 5684 8698 5740 8708
rect 7028 8764 7084 8774
rect 7028 8596 7084 8708
rect 5460 8540 5516 8596
rect 5460 8474 5516 8484
rect 5572 8540 5628 8550
rect 5124 8428 5180 8438
rect 5124 7868 5180 8372
rect 5460 8316 5516 8326
rect 5460 8204 5516 8260
rect 5460 8138 5516 8148
rect 5572 7980 5628 8484
rect 5796 8540 5852 8550
rect 5796 8316 5852 8484
rect 5796 8250 5852 8260
rect 5908 8540 5964 8550
rect 6916 8540 6972 8550
rect 6804 8484 6916 8540
rect 5908 8204 5964 8484
rect 5908 8138 5964 8148
rect 5572 7914 5628 7924
rect 3892 6794 3948 6804
rect 4228 7644 4284 7654
rect 3780 6524 3836 6534
rect 3668 4732 3724 4742
rect 3668 4284 3724 4676
rect 3780 4620 3836 6468
rect 3892 6320 3948 6330
rect 3892 6076 3948 6264
rect 3892 5648 3948 6020
rect 4228 6188 4284 7588
rect 4452 6422 4508 7700
rect 4676 7756 4732 7766
rect 4676 7532 4732 7700
rect 4788 7756 4844 7766
rect 5124 7756 5180 7812
rect 4844 7700 4956 7756
rect 4788 7690 4844 7700
rect 5124 7690 5180 7700
rect 5796 7756 5852 7766
rect 5796 7654 5852 7700
rect 5791 7644 5852 7654
rect 5847 7588 5852 7644
rect 5908 7756 5964 7766
rect 6916 7761 6972 8484
rect 7252 8540 7308 8652
rect 7252 8474 7308 8484
rect 7364 8540 7420 8550
rect 7364 8418 7420 8484
rect 7588 8540 7644 8550
rect 7252 8362 7420 8418
rect 7476 8428 7532 8438
rect 7252 8316 7308 8362
rect 7252 8250 7308 8260
rect 7252 7868 7308 7878
rect 6906 7705 6916 7761
rect 6972 7705 6982 7761
rect 5908 7654 5964 7700
rect 5908 7644 5984 7654
rect 5908 7588 5928 7644
rect 5791 7578 5847 7588
rect 5908 7578 5984 7588
rect 6916 7639 6972 7649
rect 4676 7466 4732 7476
rect 5908 7420 5964 7578
rect 6916 7471 6972 7583
rect 5796 7364 5964 7420
rect 5124 6860 5180 6870
rect 5796 6860 5852 7364
rect 5992 7196 6044 7252
rect 6100 7196 6200 7252
rect 6256 7196 6356 7252
rect 6412 7196 6512 7252
rect 6568 7196 6668 7252
rect 6724 7196 6776 7252
rect 4676 6748 4732 6758
rect 5124 6748 5180 6804
rect 4732 6692 4844 6748
rect 4676 6682 4732 6692
rect 5124 6682 5180 6692
rect 5236 6748 5292 6860
rect 5796 6794 5852 6804
rect 6132 6860 6188 6870
rect 5236 6682 5292 6692
rect 5460 6748 5516 6758
rect 4412 6361 4508 6422
rect 4564 6524 4620 6534
rect 4412 6198 4468 6361
rect 4412 6132 4468 6142
rect 3892 5582 3948 5592
rect 4004 5964 4060 5974
rect 3780 4554 3836 4564
rect 3892 5511 3948 5521
rect 3892 4956 3948 5455
rect 4004 5068 4060 5908
rect 4004 5002 4060 5012
rect 4116 5068 4172 5078
rect 3668 4218 3724 4228
rect 3780 4172 3836 4182
rect 3780 3948 3836 4116
rect 3892 4172 3948 4900
rect 3892 4106 3948 4116
rect 4004 4508 4060 4518
rect 3780 3164 3836 3892
rect 3780 3098 3836 3108
rect 3892 3164 3948 3174
rect 3556 2762 3612 2772
rect 3892 2940 3948 3108
rect 3892 2492 3948 2884
rect 3892 2426 3948 2436
rect 2772 1372 2828 1382
rect 2660 1316 2772 1372
rect 2772 1306 2828 1316
rect 3108 924 3164 2324
rect 3668 2156 3724 2166
rect 3668 1708 3724 2100
rect 3556 1596 3612 1606
rect 3444 1540 3556 1596
rect 3556 1530 3612 1540
rect 3668 1484 3724 1652
rect 3668 1372 3724 1428
rect 3668 1306 3724 1316
rect 4004 1484 4060 4452
rect 4116 4401 4172 5012
rect 4116 4335 4172 4345
rect 4228 4396 4284 6132
rect 4564 6116 4620 6468
rect 4900 6524 4956 6534
rect 4900 6300 4956 6468
rect 4900 6234 4956 6244
rect 5460 6300 5516 6692
rect 5460 6234 5516 6244
rect 5684 6748 5740 6758
rect 4544 6106 4620 6116
rect 4600 6050 4620 6106
rect 4798 6188 4854 6198
rect 4681 6076 4737 6086
rect 4544 6040 4620 6050
rect 4564 6030 4620 6040
rect 4676 6020 4681 6076
rect 4676 6010 4737 6020
rect 4452 5964 4508 5974
rect 4452 5852 4508 5908
rect 4452 5786 4508 5796
rect 4564 5959 4620 5969
rect 4452 5696 4508 5706
rect 4228 4330 4284 4340
rect 4340 5292 4396 5302
rect 4116 4264 4172 4274
rect 4116 4172 4172 4208
rect 4116 4106 4172 4116
rect 4340 4172 4396 5236
rect 4452 4396 4508 5640
rect 4564 5068 4620 5903
rect 4676 5852 4732 6010
rect 4798 5950 4854 6132
rect 5572 6188 5628 6198
rect 5236 6076 5292 6086
rect 4676 5078 4732 5796
rect 4788 5899 4854 5950
rect 5007 5964 5068 5974
rect 5236 5964 5292 6020
rect 5348 5964 5404 5974
rect 5236 5908 5348 5964
rect 4788 5701 4844 5899
rect 5007 5898 5068 5908
rect 5348 5898 5404 5908
rect 4788 5635 4844 5645
rect 4900 5852 4956 5862
rect 4676 5012 4732 5022
rect 4788 5384 4844 5394
rect 4564 5002 4620 5012
rect 4676 4951 4732 4956
rect 4671 4946 4732 4951
rect 4671 4890 4676 4946
rect 4671 4801 4732 4890
rect 4452 4330 4508 4340
rect 4340 4106 4396 4116
rect 4564 4172 4620 4284
rect 4564 4106 4620 4116
rect 4452 4060 4508 4070
rect 4116 3388 4172 3398
rect 4116 3164 4172 3332
rect 4452 3393 4508 4004
rect 4452 3327 4508 3337
rect 4564 3500 4620 3510
rect 4116 3098 4172 3108
rect 4228 3164 4284 3174
rect 4228 3052 4284 3108
rect 4564 3164 4620 3444
rect 4564 3098 4620 3108
rect 4228 2986 4284 2996
rect 4228 2828 4284 2838
rect 4228 2604 4284 2772
rect 4228 2538 4284 2548
rect 4452 2775 4508 2785
rect 4452 2380 4508 2719
rect 4676 2775 4732 4801
rect 4788 4284 4844 5328
rect 4900 5068 4956 5796
rect 5012 5292 5068 5898
rect 5572 5852 5628 6132
rect 5684 6076 5740 6692
rect 6020 6636 6076 6646
rect 6020 6188 6076 6580
rect 6132 6524 6188 6804
rect 6132 6458 6188 6468
rect 6916 6524 6972 6534
rect 6020 6122 6076 6132
rect 6916 6188 6972 6468
rect 6916 6122 6972 6132
rect 5684 6010 5740 6020
rect 5572 5786 5628 5796
rect 5796 5964 5852 5974
rect 5796 5729 5852 5908
rect 5012 5226 5068 5236
rect 5124 5673 5852 5729
rect 6916 5964 6972 5974
rect 5124 5180 5180 5673
rect 5992 5404 6044 5460
rect 6100 5404 6200 5460
rect 6256 5404 6356 5460
rect 6412 5404 6512 5460
rect 6568 5404 6668 5460
rect 6724 5404 6776 5460
rect 6132 5292 6188 5302
rect 5124 5114 5180 5124
rect 5572 5180 5628 5190
rect 4900 4508 4956 5012
rect 5460 4956 5516 5068
rect 5460 4890 5516 4900
rect 5572 4956 5628 5124
rect 5572 4890 5628 4900
rect 5684 5068 5740 5078
rect 5684 4956 5740 5012
rect 5684 4890 5740 4900
rect 6132 4956 6188 5236
rect 6356 4956 6412 4966
rect 6132 4890 6188 4900
rect 5236 4844 5292 4854
rect 4900 4442 4956 4452
rect 5012 4834 5068 4844
rect 4788 4218 4844 4228
rect 4900 4284 4956 4294
rect 4900 4172 4956 4228
rect 4900 4106 4956 4116
rect 5012 3500 5068 4778
rect 5012 3434 5068 3444
rect 5124 4722 5180 4732
rect 5012 3164 5068 3174
rect 4788 2940 4844 2950
rect 4788 2790 4844 2884
rect 4676 2709 4732 2719
rect 4228 2156 4284 2166
rect 4228 1596 4284 2100
rect 4228 1530 4284 1540
rect 4004 1372 4060 1428
rect 4340 1372 4396 1382
rect 4228 1316 4340 1372
rect 4004 1306 4060 1316
rect 4340 1306 4396 1316
rect 3108 588 3164 868
rect 4452 812 4508 2324
rect 5012 2268 5068 3108
rect 5124 2492 5180 4666
rect 5236 4172 5292 4788
rect 5908 4844 5964 4854
rect 5908 4732 5964 4788
rect 6244 4844 6300 4956
rect 6412 4900 6524 4956
rect 6356 4890 6412 4900
rect 6244 4778 6300 4788
rect 5908 4666 5964 4676
rect 6916 4284 6972 5908
rect 6916 4218 6972 4228
rect 7140 5964 7196 5974
rect 5236 4106 5292 4116
rect 5684 4172 5740 4182
rect 5236 3388 5292 3398
rect 5236 3164 5292 3332
rect 5236 3098 5292 3108
rect 5460 3164 5516 3174
rect 5460 3052 5516 3108
rect 5460 2986 5516 2996
rect 5124 2426 5180 2436
rect 5572 2380 5628 2390
rect 4676 2156 4732 2166
rect 4732 2100 4844 2156
rect 4676 2090 4732 2100
rect 4452 746 4508 756
rect 4900 1484 4956 1494
rect 4676 700 4732 710
rect 3108 522 3164 532
rect 3892 588 3948 598
rect 3892 476 3948 532
rect 4676 588 4732 644
rect 4676 522 4732 532
rect 4900 588 4956 1428
rect 5012 1372 5068 2212
rect 5124 2268 5180 2278
rect 5124 1596 5180 2212
rect 5348 2156 5404 2166
rect 5348 1988 5404 2100
rect 5124 1530 5180 1540
rect 5572 1596 5628 2324
rect 5572 1530 5628 1540
rect 5012 1306 5068 1316
rect 5684 1372 5740 4116
rect 5992 3612 6044 3668
rect 6100 3612 6200 3668
rect 6256 3612 6356 3668
rect 6412 3612 6512 3668
rect 6568 3612 6668 3668
rect 6724 3612 6776 3668
rect 5796 3388 5852 3500
rect 5796 3322 5852 3332
rect 6244 2268 6300 2278
rect 6132 2212 6244 2268
rect 6244 2202 6300 2212
rect 5992 1820 6044 1876
rect 6100 1820 6200 1876
rect 6256 1820 6356 1876
rect 6412 1820 6512 1876
rect 6568 1820 6668 1876
rect 6724 1820 6776 1876
rect 5684 700 5740 1316
rect 6020 1484 6076 1494
rect 6020 1372 6076 1428
rect 6020 1306 6076 1316
rect 6356 1372 6412 1484
rect 6356 1306 6412 1316
rect 7140 1372 7196 5908
rect 7252 5964 7308 7812
rect 7364 7868 7420 7878
rect 7364 7756 7420 7812
rect 7364 7690 7420 7700
rect 7364 7527 7420 7537
rect 7364 7420 7420 7471
rect 7364 7354 7420 7364
rect 7476 6325 7532 8372
rect 7588 8011 7644 8484
rect 7700 8540 7756 8550
rect 7700 8159 7756 8484
rect 8036 8540 8092 8652
rect 8036 8474 8092 8484
rect 8148 8540 8204 8820
rect 8148 8474 8204 8484
rect 8596 9436 8652 9446
rect 7700 8080 7796 8159
rect 7588 7943 7664 8011
rect 7608 7766 7664 7943
rect 7588 7756 7664 7766
rect 7740 7766 7796 8080
rect 8596 7868 8652 9380
rect 9044 8540 9100 11284
rect 9156 11228 9212 11340
rect 9156 11162 9212 11172
rect 9268 9548 9324 12516
rect 9492 12460 9548 13860
rect 9716 13916 9772 16436
rect 9828 15820 9884 16543
rect 9828 15754 9884 15764
rect 9940 14924 9996 16670
rect 10276 16604 10332 16716
rect 10276 16538 10332 16548
rect 10052 16380 10108 16390
rect 10052 15260 10108 16324
rect 10052 15194 10108 15204
rect 10388 15148 10444 19348
rect 11620 19404 11676 19414
rect 11060 19180 11116 19190
rect 11060 18732 11116 19124
rect 11620 19180 11676 19348
rect 12628 19404 12684 19414
rect 12404 19292 12460 19302
rect 11620 19114 11676 19124
rect 11844 19180 11900 19190
rect 11060 18666 11116 18676
rect 11844 18732 11900 19124
rect 11844 18666 11900 18676
rect 12404 18732 12460 19236
rect 12628 19292 12684 19348
rect 12740 19404 12796 19414
rect 12740 19236 12796 19348
rect 12628 19226 12684 19236
rect 12404 18666 12460 18676
rect 11620 18508 11676 18518
rect 10948 18396 11004 18406
rect 10948 18228 11004 18340
rect 11060 17612 11116 17622
rect 10836 17388 10892 17398
rect 10836 16716 10892 17332
rect 11060 16940 11116 17556
rect 11284 17612 11340 17724
rect 11284 17546 11340 17556
rect 11060 16874 11116 16884
rect 10836 16650 10892 16660
rect 11620 16380 11676 18452
rect 12740 18508 12796 18518
rect 12292 18284 12348 18294
rect 12292 17612 12348 18228
rect 12740 17948 12796 18452
rect 12740 17882 12796 17892
rect 12292 17546 12348 17556
rect 12404 17500 12460 17510
rect 11620 16314 11676 16324
rect 12068 16380 12124 16390
rect 10724 15708 10780 15718
rect 10724 15540 10780 15652
rect 11732 15708 11788 15718
rect 11508 15596 11564 15606
rect 11564 15540 11676 15596
rect 11508 15530 11564 15540
rect 10388 15082 10444 15092
rect 9940 14858 9996 14868
rect 11732 14924 11788 15652
rect 11956 15708 12012 15718
rect 11956 15596 12012 15652
rect 11956 15530 12012 15540
rect 11844 15484 11900 15494
rect 11844 14944 11900 15428
rect 11844 14878 11900 14888
rect 9492 12394 9548 12404
rect 9604 12348 9660 12460
rect 9604 12282 9660 12292
rect 9716 12124 9772 13860
rect 10052 14812 10108 14822
rect 10052 13804 10108 14756
rect 10500 14812 10556 14822
rect 10500 14588 10556 14756
rect 11172 14700 11228 14710
rect 10500 14522 10556 14532
rect 10836 14588 10892 14598
rect 10052 13738 10108 13748
rect 10388 13916 10444 13926
rect 10612 13916 10668 13926
rect 10500 13860 10612 13916
rect 10388 13804 10444 13860
rect 10612 13850 10668 13860
rect 10388 13738 10444 13748
rect 10836 13692 10892 14532
rect 10612 13244 10668 13254
rect 10500 13132 10556 13142
rect 10052 12908 10108 12918
rect 9828 12796 9884 12806
rect 9884 12740 9996 12796
rect 9828 12730 9884 12740
rect 9716 12058 9772 12068
rect 10052 12348 10108 12852
rect 10500 12908 10556 13076
rect 10500 12842 10556 12852
rect 9268 8657 9324 9492
rect 9604 11900 9660 11910
rect 9268 8591 9324 8601
rect 9492 8652 9548 8662
rect 9380 8540 9436 8550
rect 9044 8474 9100 8484
rect 9268 8520 9324 8530
rect 9156 8428 9212 8438
rect 8596 7802 8652 7812
rect 7740 7756 7801 7766
rect 7740 7700 7745 7756
rect 7588 7690 7664 7700
rect 7745 7690 7801 7700
rect 8036 7756 8092 7766
rect 7700 6860 7756 6870
rect 7700 6692 7756 6804
rect 7812 6748 7868 6758
rect 7466 6269 7476 6325
rect 7532 6269 7542 6325
rect 7476 6193 7532 6198
rect 7364 6188 7532 6193
rect 7364 6137 7476 6188
rect 7476 6122 7532 6132
rect 7252 5898 7308 5908
rect 7364 6071 7420 6081
rect 7364 5740 7420 6015
rect 7364 5674 7420 5684
rect 7588 5964 7644 5974
rect 7588 5292 7644 5908
rect 7588 5226 7644 5236
rect 7812 5292 7868 6692
rect 7812 5226 7868 5236
rect 8036 6524 8092 7700
rect 9044 7756 9100 7868
rect 9044 7690 9100 7700
rect 9156 7756 9212 8372
rect 9268 8316 9324 8464
rect 9380 8372 9436 8484
rect 9268 8260 9436 8316
rect 9380 7980 9436 8260
rect 9380 7914 9436 7924
rect 9156 7690 9212 7700
rect 9492 7756 9548 8596
rect 9604 8652 9660 11844
rect 9716 10556 9772 10566
rect 9716 10444 9772 10500
rect 9940 10444 9996 10454
rect 9716 10378 9772 10388
rect 9828 10388 9940 10444
rect 9828 9548 9884 10388
rect 9940 10378 9996 10388
rect 9828 8764 9884 9492
rect 9828 8698 9884 8708
rect 9940 10108 9996 10118
rect 9940 9436 9996 10052
rect 9604 8586 9660 8596
rect 9492 7690 9548 7700
rect 9716 8316 9772 8326
rect 8260 7532 8316 7542
rect 8260 6748 8316 7476
rect 8708 7532 8764 7542
rect 8260 6682 8316 6692
rect 8596 6860 8652 6870
rect 8036 6076 8092 6468
rect 8036 5185 8092 6020
rect 8036 5119 8092 5129
rect 8372 6320 8428 6330
rect 8026 5007 8036 5063
rect 8092 5007 8102 5063
rect 7252 4956 7308 4966
rect 7252 4844 7308 4900
rect 7812 4956 7868 4966
rect 7252 4778 7308 4788
rect 7476 4844 7532 4854
rect 7364 4172 7420 4182
rect 7364 4060 7420 4116
rect 7364 3994 7420 4004
rect 7364 3276 7420 3286
rect 7364 3164 7420 3220
rect 7364 3098 7420 3108
rect 7476 3164 7532 4788
rect 7588 4060 7644 4070
rect 7644 4004 7756 4060
rect 7588 3994 7644 4004
rect 7476 3098 7532 3108
rect 7700 3164 7756 3174
rect 7812 3164 7868 4900
rect 8036 4956 8092 5007
rect 8036 4890 8092 4900
rect 8372 4956 8428 6264
rect 8596 5852 8652 6804
rect 8596 5786 8652 5796
rect 8596 5292 8652 5302
rect 8372 4890 8428 4900
rect 8484 4956 8540 4966
rect 8484 4732 8540 4900
rect 8596 4956 8652 5236
rect 8596 4890 8652 4900
rect 8484 3836 8540 4676
rect 8484 3770 8540 3780
rect 8708 4172 8764 7476
rect 9380 6860 9436 6870
rect 9156 5852 9212 5862
rect 9156 5740 9212 5796
rect 9380 5852 9436 6804
rect 9492 6748 9548 6860
rect 9492 6682 9548 6692
rect 9380 5786 9436 5796
rect 9156 5674 9212 5684
rect 9156 5414 9212 5424
rect 8932 5292 8988 5302
rect 8260 3500 8316 3510
rect 8036 3388 8092 3398
rect 7756 3108 7868 3164
rect 7924 3164 7980 3276
rect 7700 3098 7756 3108
rect 7924 3098 7980 3108
rect 8036 3164 8092 3332
rect 8260 3276 8316 3444
rect 8708 3398 8764 4116
rect 8820 4732 8876 4742
rect 8820 4172 8876 4676
rect 8820 4106 8876 4116
rect 8708 3332 8764 3342
rect 8820 3836 8876 3846
rect 8260 3210 8316 3220
rect 8036 3098 8092 3108
rect 8708 3164 8764 3276
rect 8708 3098 8764 3108
rect 8820 3164 8876 3780
rect 8596 3052 8652 3062
rect 7476 3027 7532 3037
rect 7476 2604 7532 2971
rect 7476 2538 7532 2548
rect 7700 2940 7756 2950
rect 7140 1306 7196 1316
rect 7364 2492 7420 2502
rect 7700 2497 7756 2884
rect 8260 2940 8316 2950
rect 7690 2441 7700 2497
rect 7756 2441 7766 2497
rect 5684 634 5740 644
rect 4900 522 4956 532
rect 1932 420 2044 476
rect 1876 410 1932 420
rect 3892 410 3948 420
rect 7364 476 7420 2436
rect 7700 2375 7756 2385
rect 7588 2319 7700 2375
rect 7700 2309 7756 2319
rect 8260 2273 8316 2884
rect 8596 2716 8652 2996
rect 7588 2253 7644 2263
rect 8036 2258 8092 2268
rect 7924 2202 8036 2258
rect 8260 2207 8316 2217
rect 8484 2660 8652 2716
rect 7588 1484 7644 2197
rect 8036 2192 8092 2202
rect 8250 2095 8260 2151
rect 8316 2095 8326 2151
rect 7700 1596 7756 1708
rect 7700 1530 7756 1540
rect 7588 1418 7644 1428
rect 8148 1372 8204 1382
rect 8036 1316 8148 1372
rect 8148 1306 8204 1316
rect 8260 1036 8316 2095
rect 8484 1596 8540 2660
rect 8708 2492 8764 2502
rect 8484 1530 8540 1540
rect 8596 2380 8652 2492
rect 8596 1484 8652 2324
rect 8708 2380 8764 2436
rect 8708 2314 8764 2324
rect 8820 2380 8876 3108
rect 8820 2314 8876 2324
rect 8932 3276 8988 5236
rect 9156 4956 9212 5358
rect 9716 5297 9772 8260
rect 9716 5231 9772 5241
rect 9156 4890 9212 4900
rect 9604 5048 9660 5180
rect 9604 4060 9660 4992
rect 9604 3994 9660 4004
rect 9716 5160 9772 5170
rect 8932 2380 8988 3220
rect 9268 2604 9324 2614
rect 9268 2522 9324 2548
rect 8932 2314 8988 2324
rect 9156 2466 9324 2522
rect 9156 2380 9212 2466
rect 9156 2314 9212 2324
rect 9268 2380 9324 2390
rect 9268 2268 9324 2324
rect 9268 2202 9324 2212
rect 9604 2380 9660 2390
rect 9604 2156 9660 2324
rect 9716 2380 9772 5104
rect 9940 4396 9996 9380
rect 10052 9436 10108 12292
rect 10052 9370 10108 9380
rect 10164 12124 10220 12134
rect 10164 11340 10220 12068
rect 10164 10332 10220 11284
rect 10164 9660 10220 10276
rect 9940 4330 9996 4340
rect 10052 7644 10108 7654
rect 10052 4070 10108 7588
rect 10164 7644 10220 9604
rect 10612 9996 10668 13188
rect 10724 12908 10780 12918
rect 10724 12236 10780 12852
rect 10836 12796 10892 13636
rect 11172 13020 11228 14644
rect 11732 14028 11788 14868
rect 11732 13962 11788 13972
rect 11844 14807 11900 14817
rect 11844 13356 11900 14751
rect 11844 13290 11900 13300
rect 12068 13916 12124 16324
rect 12404 15708 12460 17444
rect 12740 16604 12796 16614
rect 12404 15642 12460 15652
rect 12516 16044 12572 16054
rect 12068 13244 12124 13860
rect 12068 13178 12124 13188
rect 11620 13132 11676 13142
rect 11620 12964 11676 13076
rect 12180 13020 12236 13030
rect 12068 12964 12180 13020
rect 11172 12954 11228 12964
rect 12180 12954 12236 12964
rect 10836 12730 10892 12740
rect 11956 12796 12012 12806
rect 11956 12460 12012 12740
rect 10724 12170 10780 12180
rect 11284 12236 11340 12246
rect 10612 9548 10668 9940
rect 10612 7756 10668 9492
rect 10724 11788 10780 11798
rect 10724 9212 10780 11732
rect 11284 11228 11340 12180
rect 11508 12236 11564 12348
rect 11508 12170 11564 12180
rect 11956 11788 12012 12404
rect 11956 11722 12012 11732
rect 11060 10332 11116 10342
rect 10948 10276 11060 10332
rect 11060 10266 11116 10276
rect 10948 9436 11004 9446
rect 10836 9380 10948 9436
rect 10948 9370 11004 9380
rect 10724 9146 10780 9156
rect 11284 8764 11340 11172
rect 11508 11228 11564 11238
rect 11732 11228 11788 11238
rect 11620 11172 11732 11228
rect 11508 11116 11564 11172
rect 11732 11162 11788 11172
rect 11508 11050 11564 11060
rect 11732 10556 11788 10566
rect 11620 10444 11676 10556
rect 11732 10412 11788 10500
rect 12404 10444 12460 10556
rect 11620 10378 11676 10388
rect 12404 10378 12460 10388
rect 11732 10332 11788 10342
rect 11956 10332 12012 10342
rect 11844 10276 11956 10332
rect 11732 9772 11788 10276
rect 11956 10266 12012 10276
rect 11732 9706 11788 9716
rect 11844 10200 11900 10210
rect 11844 9772 11900 10144
rect 11844 9706 11900 9716
rect 11508 9548 11564 9558
rect 11508 9436 11564 9492
rect 12180 9548 12236 9558
rect 12236 9492 12348 9548
rect 12180 9482 12236 9492
rect 11508 9370 11564 9380
rect 11060 8652 11116 8764
rect 11060 8586 11116 8596
rect 11284 8652 11340 8708
rect 11284 8586 11340 8596
rect 11956 8764 12012 8774
rect 10612 7690 10668 7700
rect 10164 6748 10220 7588
rect 11732 7644 11788 7654
rect 11732 7196 11788 7588
rect 11732 7130 11788 7140
rect 11956 7644 12012 8708
rect 10612 6860 10668 6870
rect 10836 6860 10892 6870
rect 10668 6804 10780 6860
rect 10612 6794 10668 6804
rect 10164 6682 10220 6692
rect 10500 6748 10556 6758
rect 10500 5964 10556 6692
rect 10836 6636 10892 6804
rect 10836 6570 10892 6580
rect 11732 6860 11788 6870
rect 10500 5898 10556 5908
rect 11284 5852 11340 5862
rect 10164 5740 10220 5750
rect 10164 5180 10220 5684
rect 10164 5114 10220 5124
rect 11284 5740 11340 5796
rect 10836 5068 10892 5078
rect 10836 4956 10892 5012
rect 11284 5068 11340 5684
rect 11396 5292 11452 5404
rect 11396 5226 11452 5236
rect 11284 5002 11340 5012
rect 10836 4890 10892 4900
rect 11620 4732 11676 4742
rect 10047 4060 10108 4070
rect 10103 4004 10108 4060
rect 10047 3994 10108 4004
rect 10052 3393 10108 3994
rect 10836 4396 10892 4406
rect 10052 3327 10108 3337
rect 10276 3388 10332 3398
rect 10276 3276 10332 3332
rect 10042 3215 10052 3271
rect 10108 3215 10220 3271
rect 10276 3210 10332 3220
rect 10388 3052 10444 3062
rect 9716 2314 9772 2324
rect 9940 2604 9996 2614
rect 9940 2380 9996 2548
rect 10388 2492 10444 2996
rect 10388 2426 10444 2436
rect 9940 2314 9996 2324
rect 10164 2380 10220 2390
rect 9604 2090 9660 2100
rect 10164 2156 10220 2324
rect 10164 2090 10220 2100
rect 10500 2380 10556 2390
rect 10500 2268 10556 2324
rect 10836 2380 10892 4340
rect 11508 4060 11564 4070
rect 11620 4060 11676 4676
rect 11564 4004 11676 4060
rect 11732 4060 11788 6804
rect 11956 6865 12012 7588
rect 12516 8540 12572 15988
rect 12740 15932 12796 16548
rect 12852 16604 12908 19908
rect 12964 18284 13020 18294
rect 12964 17836 13020 18228
rect 12964 17770 13020 17780
rect 13076 17276 13132 20132
rect 13636 20188 13692 20198
rect 13636 20076 13692 20132
rect 13300 19964 13356 19974
rect 13188 19908 13300 19964
rect 13300 19898 13356 19908
rect 13300 17388 13356 17398
rect 13356 17332 13468 17388
rect 13300 17322 13356 17332
rect 13076 17210 13132 17220
rect 13524 16828 13580 16838
rect 12852 16538 12908 16548
rect 12964 16604 13020 16614
rect 12740 15866 12796 15876
rect 12964 14924 13020 16548
rect 13524 15820 13580 16772
rect 13524 15754 13580 15764
rect 12964 14812 13020 14868
rect 12964 14746 13020 14756
rect 13076 15708 13132 15718
rect 13076 14680 13132 15652
rect 12964 14624 13132 14680
rect 13188 14812 13244 14822
rect 13188 14644 13244 14756
rect 12740 14028 12796 14140
rect 12740 13962 12796 13972
rect 12852 13804 12908 13814
rect 12740 13132 12796 13244
rect 12740 13066 12796 13076
rect 12628 12908 12684 12918
rect 12628 12348 12684 12852
rect 12628 12282 12684 12292
rect 12740 12796 12796 12806
rect 12628 11228 12684 11238
rect 12628 9436 12684 11172
rect 12740 11004 12796 12740
rect 12852 12236 12908 13748
rect 12964 13356 13020 14624
rect 13300 14028 13356 14038
rect 13300 13916 13356 13972
rect 13300 13850 13356 13860
rect 13636 13580 13692 20020
rect 14084 18732 14140 20244
rect 14308 20300 14364 20412
rect 14308 20234 14364 20244
rect 16772 20300 16828 20310
rect 14084 18666 14140 18676
rect 14868 20188 14924 20198
rect 14532 18508 14588 18620
rect 14532 18442 14588 18452
rect 14756 18508 14812 18518
rect 13748 18396 13804 18406
rect 13748 16176 13804 18340
rect 14420 18396 14476 18406
rect 14308 18172 14364 18182
rect 14308 17276 14364 18116
rect 14084 16716 14140 16726
rect 13748 16120 13916 16176
rect 13636 13514 13692 13524
rect 13748 16044 13804 16054
rect 12964 13290 13020 13300
rect 12852 12170 12908 12180
rect 13412 12908 13468 12918
rect 13412 12348 13468 12852
rect 13748 12796 13804 15988
rect 13860 15148 13916 16120
rect 13860 15082 13916 15092
rect 14084 14028 14140 16660
rect 14308 15036 14364 17220
rect 14420 16828 14476 18340
rect 14756 18284 14812 18452
rect 14868 18396 14924 20132
rect 16772 20188 16828 20244
rect 18116 20300 18172 20310
rect 16772 20122 16828 20132
rect 16996 20188 17052 20198
rect 15428 19404 15484 19414
rect 15316 19348 15428 19404
rect 15316 18732 15372 19348
rect 15428 19338 15484 19348
rect 15652 19404 15708 19414
rect 15316 18666 15372 18676
rect 15652 19292 15708 19348
rect 16996 19404 17052 20132
rect 15092 18508 15148 18518
rect 14980 18452 15092 18508
rect 15092 18442 15148 18452
rect 14868 18340 15036 18396
rect 14756 18218 14812 18228
rect 14756 17500 14812 17510
rect 14756 16940 14812 17444
rect 14756 16874 14812 16884
rect 14644 16828 14700 16838
rect 14532 16772 14644 16828
rect 14420 16762 14476 16772
rect 14644 16762 14700 16772
rect 14980 16716 15036 18340
rect 14308 14970 14364 14980
rect 14644 15596 14700 15606
rect 14644 14924 14700 15540
rect 14532 14700 14588 14710
rect 14532 14145 14588 14644
rect 14532 14079 14588 14089
rect 14644 14023 14700 14868
rect 14084 13132 14140 13972
rect 14522 13967 14532 14023
rect 14588 13967 14700 14023
rect 14084 13066 14140 13076
rect 14644 13020 14700 13967
rect 14644 12954 14700 12964
rect 14756 14028 14812 14038
rect 13524 12460 13580 12572
rect 13524 12394 13580 12404
rect 13748 12460 13804 12740
rect 13748 12394 13804 12404
rect 14756 12348 14812 13972
rect 14980 12908 15036 16660
rect 14980 12842 15036 12852
rect 15092 17948 15148 17958
rect 15092 15708 15148 17892
rect 15428 17612 15484 17622
rect 15428 17500 15484 17556
rect 15652 17612 15708 19236
rect 16772 19292 16828 19302
rect 16772 19180 16828 19236
rect 16996 19292 17052 19348
rect 16996 19226 17052 19236
rect 17444 19292 17500 19302
rect 16772 19114 16828 19124
rect 17332 19180 17388 19190
rect 16408 18844 16460 18900
rect 16516 18844 16616 18900
rect 16672 18844 16772 18900
rect 16828 18844 16928 18900
rect 16984 18844 17084 18900
rect 17140 18844 17192 18900
rect 15652 17546 15708 17556
rect 16548 18732 16604 18742
rect 16548 18396 16604 18676
rect 15428 17434 15484 17444
rect 16100 17276 16156 17286
rect 15540 16716 15596 16726
rect 15540 16604 15596 16660
rect 15540 16538 15596 16548
rect 15652 16604 15708 16614
rect 15092 12572 15148 15652
rect 15652 16380 15708 16548
rect 15316 13020 15372 13132
rect 15316 12954 15372 12964
rect 15540 13020 15596 13030
rect 15540 12852 15596 12964
rect 14868 12460 14924 12572
rect 15092 12506 15148 12516
rect 15316 12572 15372 12582
rect 14868 12394 14924 12404
rect 13412 12236 13468 12292
rect 13412 12170 13468 12180
rect 14084 12236 14140 12348
rect 14756 12282 14812 12292
rect 15092 12236 15148 12246
rect 14980 12180 15092 12236
rect 14084 12170 14140 12180
rect 15092 12170 15148 12180
rect 12964 12124 13020 12134
rect 12964 12012 13020 12068
rect 12964 11946 13020 11956
rect 13860 12124 13916 12134
rect 12852 11340 12908 11452
rect 13748 11340 13804 11350
rect 12852 11274 12908 11284
rect 13412 11228 13468 11340
rect 13412 11162 13468 11172
rect 13524 11116 13580 11228
rect 13524 11050 13580 11060
rect 12740 10668 12796 10948
rect 13748 10892 13804 11284
rect 13748 10826 13804 10836
rect 12740 10602 12796 10612
rect 13412 10668 13468 10678
rect 12964 9548 13020 9558
rect 13020 9492 13132 9548
rect 12964 9482 13020 9492
rect 12628 9370 12684 9380
rect 12740 9212 12796 9222
rect 12628 9156 12740 9212
rect 12740 9146 12796 9156
rect 13188 9212 13244 9222
rect 12516 7084 12572 8484
rect 13076 7756 13132 7766
rect 13076 7644 13132 7700
rect 13076 7578 13132 7588
rect 12516 7018 12572 7028
rect 12740 7196 12796 7206
rect 12740 6972 12796 7140
rect 12964 7196 13020 7206
rect 11956 6799 12012 6809
rect 12516 6870 12572 6960
rect 12740 6906 12796 6916
rect 12852 7084 12908 7094
rect 12516 6804 12572 6814
rect 12628 6748 12684 6758
rect 11946 6687 11956 6743
rect 12012 6687 12124 6743
rect 12516 6692 12628 6748
rect 12516 6524 12572 6692
rect 12628 6682 12684 6692
rect 12516 6458 12572 6468
rect 12404 5964 12460 5974
rect 12180 5857 12236 5867
rect 11956 4956 12012 4966
rect 11956 4844 12012 4900
rect 11956 4778 12012 4788
rect 11508 3994 11564 4004
rect 11732 3994 11788 4004
rect 11508 3164 11564 3276
rect 11508 3098 11564 3108
rect 12180 2604 12236 5801
rect 12404 5628 12460 5908
rect 12516 5969 12572 5979
rect 12572 5913 12684 5969
rect 12516 5903 12572 5913
rect 12740 5857 12796 5867
rect 12628 5801 12740 5857
rect 12740 5791 12796 5801
rect 12404 5562 12460 5572
rect 12628 5735 12684 5745
rect 12628 5292 12684 5679
rect 12628 5226 12684 5236
rect 12740 5628 12796 5638
rect 12740 5180 12796 5572
rect 12404 5068 12460 5078
rect 12404 4396 12460 5012
rect 12404 4330 12460 4340
rect 12740 4172 12796 5124
rect 12740 4106 12796 4116
rect 12852 4172 12908 7028
rect 12964 6748 13020 7140
rect 13188 7084 13244 9156
rect 13412 9212 13468 10612
rect 13636 10444 13692 10454
rect 13524 10388 13636 10444
rect 13636 10378 13692 10388
rect 13748 9548 13804 9660
rect 13748 9482 13804 9492
rect 13412 9146 13468 9156
rect 13636 9436 13692 9446
rect 13636 8764 13692 9380
rect 13860 9314 13916 12068
rect 14420 12124 14476 12134
rect 14420 11956 14476 12068
rect 14756 12124 14812 12134
rect 14532 12012 14588 12022
rect 14196 11228 14252 11238
rect 14196 11060 14252 11172
rect 14420 11004 14476 11014
rect 14308 10948 14420 11004
rect 14420 10938 14476 10948
rect 14298 10831 14308 10887
rect 14364 10831 14374 10887
rect 14196 10556 14252 10566
rect 14196 10332 14252 10500
rect 14308 10444 14364 10831
rect 14532 10556 14588 11956
rect 14532 10490 14588 10500
rect 14308 10378 14364 10388
rect 14196 10266 14252 10276
rect 14084 10108 14140 10118
rect 13972 9548 14028 9558
rect 13972 9426 14028 9492
rect 14084 9548 14140 10052
rect 14756 9772 14812 12068
rect 14868 10444 14924 10454
rect 14868 10276 14924 10388
rect 15092 10332 15148 10342
rect 14756 9706 14812 9716
rect 14980 9772 15036 9782
rect 14980 9670 15036 9716
rect 14868 9614 15036 9670
rect 14084 9482 14140 9492
rect 14196 9548 14252 9558
rect 14196 9436 14252 9492
rect 13972 9370 14140 9426
rect 14196 9370 14252 9380
rect 14420 9548 14476 9558
rect 14532 9548 14588 9558
rect 14476 9492 14532 9548
rect 13860 9258 14028 9314
rect 13636 8698 13692 8708
rect 13300 8652 13356 8662
rect 13300 7756 13356 8596
rect 13300 7690 13356 7700
rect 13412 7980 13468 7990
rect 13188 7018 13244 7028
rect 13300 6860 13356 6870
rect 13188 6804 13300 6860
rect 13300 6794 13356 6804
rect 12964 6682 13020 6692
rect 12964 5969 13020 5979
rect 12964 5852 13020 5913
rect 12964 5628 13020 5796
rect 12964 5562 13020 5572
rect 13300 5852 13356 5862
rect 12964 4956 13020 4966
rect 13020 4900 13132 4956
rect 12964 4890 13020 4900
rect 12516 3276 12572 3286
rect 12572 3220 12684 3276
rect 12516 3210 12572 3220
rect 12852 3174 12908 4116
rect 13300 4396 13356 5796
rect 13412 4961 13468 7924
rect 13636 7532 13692 7542
rect 13636 6860 13692 7476
rect 13636 6794 13692 6804
rect 13860 6972 13916 6982
rect 13860 6748 13916 6916
rect 13972 6860 14028 9258
rect 14084 7308 14140 9370
rect 14084 7242 14140 7252
rect 14196 8876 14252 8886
rect 13972 6794 14028 6804
rect 13860 6682 13916 6692
rect 14196 6604 14252 8820
rect 14420 8540 14476 9492
rect 14532 9482 14588 9492
rect 14644 9548 14700 9558
rect 14420 7980 14476 8484
rect 14420 7914 14476 7924
rect 14532 9304 14588 9314
rect 14532 7756 14588 9248
rect 14644 8988 14700 9492
rect 14868 9553 14924 9614
rect 14868 9487 14924 9497
rect 14980 9548 15036 9558
rect 14644 8922 14700 8932
rect 14868 9416 14924 9426
rect 14644 8540 14700 8550
rect 14644 8428 14700 8484
rect 14756 8540 14812 8652
rect 14756 8474 14812 8484
rect 14644 8362 14700 8372
rect 14868 8428 14924 9360
rect 14756 7980 14812 7990
rect 14756 7812 14812 7924
rect 14186 6542 14252 6604
rect 14308 6636 14364 6646
rect 14186 6086 14242 6542
rect 14176 6030 14186 6086
rect 14242 6030 14252 6086
rect 13636 5964 13692 5974
rect 13692 5908 13804 5964
rect 14196 5959 14252 5969
rect 13636 5898 13692 5908
rect 13524 5740 13580 5750
rect 13524 5078 13580 5684
rect 13524 5012 13580 5022
rect 13412 4895 13468 4905
rect 13636 4956 13692 4966
rect 13860 4956 13916 4966
rect 13692 4900 13804 4956
rect 13636 4890 13692 4900
rect 13300 3388 13356 4340
rect 13412 4824 13468 4834
rect 13412 4396 13468 4768
rect 13412 4330 13468 4340
rect 13860 4284 13916 4900
rect 13300 3322 13356 3332
rect 13636 3500 13692 3510
rect 12832 3164 12908 3174
rect 12888 3108 12908 3164
rect 12964 3164 13025 3174
rect 13188 3164 13244 3174
rect 13025 3108 13132 3164
rect 12832 3098 12888 3108
rect 12964 3098 13025 3108
rect 12292 3052 12348 3062
rect 12292 2940 12348 2996
rect 12292 2874 12348 2884
rect 12964 2940 13020 3098
rect 12964 2874 13020 2884
rect 10836 2314 10892 2324
rect 11060 2380 11116 2390
rect 11732 2380 11788 2390
rect 11620 2324 11732 2380
rect 11060 2268 11116 2324
rect 11732 2314 11788 2324
rect 10388 2044 10444 2054
rect 9940 1596 9996 1606
rect 9828 1540 9940 1596
rect 9940 1530 9996 1540
rect 8596 1418 8652 1428
rect 9828 1372 9884 1382
rect 9716 1316 9828 1372
rect 9828 1306 9884 1316
rect 10388 1372 10444 1988
rect 10500 1601 10556 2212
rect 10612 2156 10668 2268
rect 11060 2202 11116 2212
rect 11172 2268 11228 2278
rect 10612 2090 10668 2100
rect 11172 2044 11228 2212
rect 11172 1978 11228 1988
rect 12068 2268 12124 2278
rect 10500 1535 10556 1545
rect 8708 1260 8764 1270
rect 8764 1204 8876 1260
rect 8708 1194 8764 1204
rect 8260 970 8316 980
rect 8708 924 8764 934
rect 8708 588 8764 868
rect 9268 700 9324 710
rect 9156 644 9268 700
rect 9268 634 9324 644
rect 10388 700 10444 1316
rect 10388 634 10444 644
rect 10500 1464 10556 1474
rect 8708 522 8764 532
rect 10500 588 10556 1408
rect 10500 522 10556 532
rect 11396 1372 11452 1382
rect 11396 588 11452 1316
rect 12068 1372 12124 2212
rect 12068 1306 12124 1316
rect 11396 522 11452 532
rect 11508 812 11564 822
rect 11508 588 11564 756
rect 12180 812 12236 2548
rect 12292 2380 12348 2390
rect 13188 2380 13244 3108
rect 12348 2324 12460 2380
rect 12292 2314 12348 2324
rect 13188 2314 13244 2324
rect 13300 2492 13356 2502
rect 13300 1596 13356 2436
rect 13524 2380 13580 2390
rect 13524 2268 13580 2324
rect 13300 1530 13356 1540
rect 13412 2212 13580 2268
rect 13412 1489 13468 2212
rect 13524 2146 13580 2156
rect 13524 1596 13580 2090
rect 13636 2044 13692 3444
rect 13860 3388 13916 4228
rect 13860 3322 13916 3332
rect 13972 4956 14028 4966
rect 13636 1978 13692 1988
rect 13524 1530 13580 1540
rect 13972 1708 14028 4900
rect 14084 3164 14140 3174
rect 14084 3052 14140 3108
rect 14196 3164 14252 5903
rect 14308 4844 14364 6580
rect 14532 6626 14588 7700
rect 14756 7196 14812 7206
rect 14756 7084 14812 7140
rect 14756 7018 14812 7028
rect 14756 6860 14812 6870
rect 14644 6804 14756 6860
rect 14644 6748 14700 6804
rect 14756 6794 14812 6804
rect 14644 6682 14700 6692
rect 14868 6636 14924 8372
rect 14980 8316 15036 9492
rect 15092 9100 15148 10276
rect 15204 10108 15260 10118
rect 15204 9682 15260 10052
rect 15204 9616 15260 9626
rect 15316 9212 15372 12516
rect 15540 12124 15596 12134
rect 15540 11956 15596 12068
rect 15652 11900 15708 16324
rect 16100 16604 16156 17220
rect 16548 17276 16604 18340
rect 17332 18508 17388 19124
rect 16884 17500 16940 17612
rect 16884 17434 16940 17444
rect 17332 17500 17388 18452
rect 17444 19180 17500 19236
rect 17444 18508 17500 19124
rect 18116 19180 18172 20244
rect 19348 20300 19404 20310
rect 18788 20188 18844 20198
rect 18788 20076 18844 20132
rect 18788 20010 18844 20020
rect 19348 19516 19404 20244
rect 20468 20300 20524 20356
rect 20468 20234 20524 20244
rect 21140 20300 21196 20412
rect 21140 20234 21196 20244
rect 19908 20188 19964 20198
rect 19348 19450 19404 19460
rect 19684 19852 19740 19862
rect 18116 19114 18172 19124
rect 18452 19404 18508 19414
rect 17561 18508 17617 18518
rect 17444 18442 17500 18452
rect 17556 18452 17561 18508
rect 17556 18442 17617 18452
rect 17332 17434 17388 17444
rect 16548 17210 16604 17220
rect 16408 17052 16460 17108
rect 16516 17052 16616 17108
rect 16672 17052 16772 17108
rect 16828 17052 16928 17108
rect 16984 17052 17084 17108
rect 17140 17052 17192 17108
rect 16884 16940 16940 16950
rect 16884 16772 16940 16884
rect 16660 16716 16716 16726
rect 16716 16660 16828 16716
rect 16660 16650 16716 16660
rect 15988 13936 16044 13946
rect 15652 11834 15708 11844
rect 15764 13916 15820 13926
rect 15876 13880 15988 13936
rect 15988 13870 16044 13880
rect 15652 11228 15708 11238
rect 15428 10556 15484 10566
rect 15484 10500 15596 10556
rect 15428 10490 15484 10500
rect 15428 10332 15484 10342
rect 15428 9558 15484 10276
rect 15652 9682 15708 11172
rect 15428 9492 15484 9502
rect 15540 9558 15596 9682
rect 15540 9492 15596 9502
rect 15652 9548 15708 9626
rect 15652 9482 15708 9492
rect 15540 9324 15596 9334
rect 15306 9156 15316 9212
rect 15372 9156 15382 9212
rect 15540 9100 15596 9268
rect 15306 9044 15316 9100
rect 15372 9044 15382 9100
rect 15092 9034 15148 9044
rect 15316 8764 15372 9044
rect 15540 9034 15596 9044
rect 15428 8988 15484 8998
rect 15428 8876 15484 8932
rect 15428 8810 15484 8820
rect 15764 8876 15820 13860
rect 15988 13799 16044 13809
rect 15876 12124 15932 12236
rect 15876 12058 15932 12068
rect 15988 11992 16044 13743
rect 15764 8810 15820 8820
rect 15876 11936 16044 11992
rect 16100 12012 16156 16548
rect 17220 15596 17276 15606
rect 17220 15428 17276 15540
rect 16408 15260 16460 15316
rect 16516 15260 16616 15316
rect 16672 15260 16772 15316
rect 16828 15260 16928 15316
rect 16984 15260 17084 15316
rect 17140 15260 17192 15316
rect 17220 14924 17276 14934
rect 16996 14812 17052 14822
rect 16212 14588 16268 14598
rect 16212 14140 16268 14532
rect 16996 14588 17052 14756
rect 17220 14812 17276 14868
rect 17220 14746 17276 14756
rect 16996 14522 17052 14532
rect 16212 14074 16268 14084
rect 16436 14364 16492 14374
rect 16436 13916 16492 14308
rect 16436 13804 16492 13860
rect 16548 13916 16604 13926
rect 16604 13860 16716 13916
rect 16548 13850 16604 13860
rect 16436 13738 16492 13748
rect 17332 13804 17388 13814
rect 17556 13804 17612 18442
rect 18452 18396 18508 19348
rect 19124 19404 19180 19414
rect 18788 19292 18844 19302
rect 18676 19236 18788 19292
rect 18788 19226 18844 19236
rect 19124 19292 19180 19348
rect 19460 19292 19516 19302
rect 19348 19236 19460 19292
rect 19124 19226 19180 19236
rect 19460 19226 19516 19236
rect 19684 19292 19740 19796
rect 19796 19292 19852 19302
rect 19684 19236 19796 19292
rect 18452 18330 18508 18340
rect 18676 18396 18732 18406
rect 17444 13748 17556 13804
rect 16408 13468 16460 13524
rect 16516 13468 16616 13524
rect 16672 13468 16772 13524
rect 16828 13468 16928 13524
rect 16984 13468 17084 13524
rect 17140 13468 17192 13524
rect 16884 13020 16940 13030
rect 16884 12348 16940 12964
rect 16884 12282 16940 12292
rect 16100 11946 16156 11956
rect 15876 10444 15932 11936
rect 16408 11676 16460 11732
rect 16516 11676 16616 11732
rect 16672 11676 16772 11732
rect 16828 11676 16928 11732
rect 16984 11676 17084 11732
rect 17140 11676 17192 11732
rect 17108 11340 17164 11350
rect 17164 11284 17276 11340
rect 17108 11274 17164 11284
rect 16212 11228 16268 11238
rect 16212 11087 16268 11172
rect 15316 8698 15372 8708
rect 15652 8652 15708 8662
rect 14980 8250 15036 8260
rect 15204 8540 15260 8550
rect 15204 7896 15260 8484
rect 15184 7844 15260 7896
rect 15428 8540 15484 8550
rect 14980 7756 15036 7766
rect 14980 7644 15036 7700
rect 14980 7578 15036 7588
rect 15184 7428 15240 7844
rect 15428 7654 15484 8484
rect 15652 8545 15708 8596
rect 15652 8479 15708 8489
rect 15764 8540 15820 8550
rect 15652 8408 15708 8418
rect 15764 8372 15820 8484
rect 15652 7980 15708 8352
rect 15652 7914 15708 7924
rect 15876 7873 15932 10388
rect 16212 11004 16268 11014
rect 16212 10444 16268 10948
rect 17332 11004 17388 13748
rect 17556 13738 17612 13748
rect 17668 17388 17724 17398
rect 17668 16716 17724 17332
rect 18676 16945 18732 18340
rect 19012 18396 19068 18406
rect 19012 17724 19068 18340
rect 19012 17658 19068 17668
rect 19572 17500 19628 17510
rect 18788 17388 18844 17500
rect 18788 17322 18844 17332
rect 19572 17388 19628 17444
rect 19572 17322 19628 17332
rect 18676 16879 18732 16889
rect 18666 16767 18676 16823
rect 18732 16767 18742 16823
rect 17556 13356 17612 13366
rect 17332 10938 17388 10948
rect 17444 13132 17500 13142
rect 17444 10556 17500 13076
rect 17556 13020 17612 13300
rect 17556 12852 17612 12964
rect 17556 12144 17612 12236
rect 17556 12078 17612 12088
rect 17444 10490 17500 10500
rect 17556 12007 17612 12017
rect 17556 10892 17612 11951
rect 16212 10378 16268 10388
rect 15988 10332 16044 10342
rect 16324 10332 16380 10342
rect 15988 10164 16044 10276
rect 16212 10276 16324 10322
rect 16212 10266 16380 10276
rect 15988 9660 16044 9772
rect 15988 9594 16044 9604
rect 16100 9436 16156 9446
rect 16100 8988 16156 9380
rect 16212 9436 16268 10266
rect 16408 9884 16460 9940
rect 16516 9884 16616 9940
rect 16672 9884 16772 9940
rect 16828 9884 16928 9940
rect 16984 9884 17084 9940
rect 17140 9884 17192 9940
rect 16212 9370 16268 9380
rect 17108 9548 17164 9558
rect 16100 8922 16156 8932
rect 16772 8988 16828 8998
rect 16324 8876 16380 8886
rect 16100 8764 16156 8774
rect 16100 8596 16156 8708
rect 16324 8764 16380 8820
rect 16324 8698 16380 8708
rect 16772 8764 16828 8932
rect 16772 8698 16828 8708
rect 15876 7807 15932 7817
rect 15988 8540 16044 8550
rect 17108 8540 17164 9492
rect 17332 9324 17388 9334
rect 17332 9100 17388 9268
rect 17556 9110 17612 10836
rect 17668 9996 17724 16660
rect 17780 16044 17836 16054
rect 17780 15820 17836 15988
rect 17780 15754 17836 15764
rect 18340 16044 18396 16054
rect 18340 14924 18396 15988
rect 18340 14028 18396 14868
rect 18340 13962 18396 13972
rect 18116 13132 18172 13142
rect 18004 12908 18060 12918
rect 17892 12852 18004 12908
rect 18004 12842 18060 12852
rect 18004 12348 18060 12358
rect 18004 12180 18060 12292
rect 18116 12124 18172 13076
rect 18564 13020 18620 13030
rect 18228 12796 18284 12806
rect 18228 12460 18284 12740
rect 18228 12394 18284 12404
rect 18116 12058 18172 12068
rect 18564 12124 18620 12964
rect 18228 11228 18284 11238
rect 18116 11172 18228 11228
rect 18228 11162 18284 11172
rect 18452 11228 18508 11238
rect 18340 10439 18396 10449
rect 17668 9930 17724 9940
rect 18228 10332 18284 10342
rect 18228 9772 18284 10276
rect 18228 9706 18284 9716
rect 17668 9436 17724 9548
rect 17668 9370 17724 9380
rect 17892 9436 17948 9446
rect 17948 9380 18060 9436
rect 17892 9370 17948 9380
rect 18004 9212 18060 9380
rect 18340 9324 18396 10383
rect 18452 9660 18508 11172
rect 18564 11004 18620 12068
rect 18564 10938 18620 10948
rect 18676 10556 18732 16767
rect 18788 16604 18844 16614
rect 18788 15820 18844 16548
rect 19348 16604 19404 16614
rect 18788 14924 18844 15764
rect 18900 15820 18956 15830
rect 18900 15652 18956 15764
rect 18844 14868 18956 14924
rect 18788 14858 18844 14868
rect 18788 14028 18844 14038
rect 18788 13804 18844 13972
rect 18788 13738 18844 13748
rect 18900 14028 18956 14868
rect 19012 14812 19068 14822
rect 19012 14364 19068 14756
rect 19012 14298 19068 14308
rect 18788 13244 18844 13254
rect 18788 13020 18844 13188
rect 18788 12954 18844 12964
rect 18900 11228 18956 13972
rect 19124 13804 19180 13814
rect 19124 13356 19180 13748
rect 19124 13290 19180 13300
rect 18900 11162 18956 11172
rect 19124 13020 19180 13030
rect 19124 12348 19180 12964
rect 19348 12684 19404 16548
rect 19460 16604 19516 16614
rect 19460 16436 19516 16548
rect 19572 13916 19628 13926
rect 19460 13356 19516 13366
rect 19460 13132 19516 13300
rect 19460 13066 19516 13076
rect 19572 13132 19628 13860
rect 19572 12796 19628 13076
rect 19684 13020 19740 19236
rect 19796 19226 19852 19236
rect 19796 18508 19852 18518
rect 19796 18172 19852 18452
rect 19796 18106 19852 18116
rect 19908 15036 19964 20132
rect 20692 19180 20748 19190
rect 20356 18732 20412 18742
rect 20356 18620 20412 18676
rect 20356 18554 20412 18564
rect 20468 18508 20524 18518
rect 20468 18396 20524 18452
rect 20468 18330 20524 18340
rect 20244 17500 20300 17510
rect 20244 17332 20300 17444
rect 20356 16716 20412 16726
rect 20356 15932 20412 16660
rect 20468 16604 20524 16614
rect 20468 16049 20524 16548
rect 20468 15983 20524 15993
rect 20356 15866 20412 15876
rect 20468 15912 20524 15922
rect 20132 15708 20188 15718
rect 20132 15148 20188 15652
rect 20132 15082 20188 15092
rect 20244 15596 20300 15606
rect 19908 14970 19964 14980
rect 19908 14028 19964 14038
rect 19964 13972 20076 14028
rect 19908 13962 19964 13972
rect 19684 12954 19740 12964
rect 20132 13132 20188 13142
rect 19572 12730 19628 12740
rect 20132 12801 20188 13076
rect 20244 13132 20300 15540
rect 20300 13076 20412 13132
rect 20244 13066 20300 13076
rect 20132 12735 20188 12745
rect 19348 12618 19404 12628
rect 20122 12623 20132 12679
rect 20188 12623 20198 12679
rect 18676 10490 18732 10500
rect 19124 10220 19180 12292
rect 20132 12348 20188 12623
rect 20132 12282 20188 12292
rect 19796 12236 19852 12246
rect 19236 12124 19292 12134
rect 19236 11956 19292 12068
rect 19796 12012 19852 12180
rect 19796 11946 19852 11956
rect 20244 12124 20300 12134
rect 20244 11340 20300 12068
rect 20468 12124 20524 15856
rect 20580 15800 20636 15810
rect 20580 13356 20636 15744
rect 20692 14476 20748 19124
rect 20804 19180 20860 19190
rect 20804 19012 20860 19124
rect 21140 18508 21196 18518
rect 21140 18340 21196 18452
rect 21364 18508 21420 20972
rect 22372 20300 22428 20310
rect 22260 20244 22372 20300
rect 22260 20188 22316 20244
rect 22372 20234 22428 20244
rect 22260 20122 22316 20132
rect 21364 18442 21420 18452
rect 21476 20076 21532 20086
rect 20916 18284 20972 18294
rect 20692 14410 20748 14420
rect 20804 17388 20860 17398
rect 20804 14252 20860 17332
rect 20916 14700 20972 18228
rect 21476 17836 21532 20020
rect 21588 19628 21644 19638
rect 21588 19292 21644 19572
rect 21588 19226 21644 19236
rect 21812 19180 21868 19190
rect 21700 18620 21756 18630
rect 21588 18564 21700 18620
rect 21700 18554 21756 18564
rect 21476 17770 21532 17780
rect 21812 18508 21868 19124
rect 21476 17500 21532 17510
rect 21364 17444 21476 17500
rect 21364 17388 21420 17444
rect 21476 17434 21532 17444
rect 21364 17322 21420 17332
rect 21812 16828 21868 18452
rect 22148 19180 22204 19190
rect 22148 17612 22204 19124
rect 22484 18508 22540 20972
rect 22708 19180 22764 20972
rect 23156 20300 23212 20310
rect 22820 20076 22876 20086
rect 22820 19745 22876 20020
rect 22820 19679 22876 19689
rect 22820 19608 22876 19618
rect 22820 19292 22876 19552
rect 22820 19226 22876 19236
rect 22708 19114 22764 19124
rect 22484 18340 22540 18452
rect 23156 18396 23212 20244
rect 22260 18284 22316 18294
rect 22260 18060 22316 18228
rect 22932 18284 22988 18396
rect 23156 18330 23212 18340
rect 23492 20076 23548 20086
rect 22932 18218 22988 18228
rect 22260 17994 22316 18004
rect 22148 17546 22204 17556
rect 22708 17500 22764 17510
rect 22596 17444 22708 17500
rect 21812 16762 21868 16772
rect 22036 17388 22092 17398
rect 21140 16604 21196 16614
rect 21140 15932 21196 16548
rect 22036 16268 22092 17332
rect 22596 17388 22652 17444
rect 22708 17434 22764 17444
rect 22596 17322 22652 17332
rect 23380 16828 23436 16838
rect 22260 16716 22316 16726
rect 22148 16660 22260 16716
rect 22148 16604 22204 16660
rect 22260 16650 22316 16660
rect 22148 16538 22204 16548
rect 22036 16202 22092 16212
rect 22708 16492 22764 16502
rect 21140 15866 21196 15876
rect 21252 15708 21308 15718
rect 21140 15652 21252 15708
rect 21140 15596 21196 15652
rect 21252 15642 21308 15652
rect 21700 15657 21812 15713
rect 21868 15657 21878 15713
rect 21140 15530 21196 15540
rect 21700 15148 21756 15657
rect 21700 15082 21756 15092
rect 21812 15591 21868 15601
rect 21140 15036 21196 15046
rect 21140 14924 21196 14980
rect 21140 14858 21196 14868
rect 20916 14634 20972 14644
rect 20804 14186 20860 14196
rect 21140 14028 21196 14038
rect 20580 13290 20636 13300
rect 20804 13804 20860 13814
rect 20804 13356 20860 13748
rect 20692 13020 20748 13030
rect 20692 12913 20748 12964
rect 20804 13020 20860 13300
rect 20804 12954 20860 12964
rect 21028 13132 21084 13142
rect 21028 13020 21084 13076
rect 21028 12954 21084 12964
rect 20692 12847 20748 12857
rect 20682 12735 20692 12791
rect 20748 12735 20758 12791
rect 20468 12012 20524 12068
rect 20468 11946 20524 11956
rect 20692 12124 20748 12735
rect 20020 11228 20076 11238
rect 19908 11116 19964 11126
rect 19908 10892 19964 11060
rect 19908 10826 19964 10836
rect 19460 10464 19516 10474
rect 19348 10352 19404 10464
rect 19348 10286 19404 10296
rect 19460 10332 19516 10408
rect 20020 10444 20076 11172
rect 20020 10378 20076 10388
rect 19460 10266 19516 10276
rect 19124 10154 19180 10164
rect 19348 10220 19404 10230
rect 18452 9594 18508 9604
rect 18340 9258 18396 9268
rect 18788 9436 18844 9446
rect 18004 9156 18172 9212
rect 17332 9034 17388 9044
rect 17546 9048 17612 9110
rect 17546 8764 17602 9048
rect 17546 8698 17602 8708
rect 17658 8988 17714 8998
rect 17658 8570 17714 8932
rect 18116 8886 18172 9156
rect 18676 9100 18732 9110
rect 17775 8876 17831 8886
rect 17912 8876 17968 8886
rect 17831 8820 17836 8876
rect 17775 8810 17836 8820
rect 17780 8652 17836 8810
rect 17892 8820 17912 8876
rect 18116 8876 18192 8886
rect 18116 8820 18136 8876
rect 17892 8810 17968 8820
rect 18136 8810 18192 8820
rect 17892 8764 17948 8810
rect 17892 8698 17948 8708
rect 17780 8586 17836 8596
rect 17098 8484 17108 8540
rect 17164 8484 17174 8540
rect 17658 8512 17724 8570
rect 15988 7756 16044 8484
rect 16324 8428 16380 8438
rect 17220 8428 17276 8438
rect 16212 8372 16324 8428
rect 17108 8372 17220 8428
rect 15876 7736 15932 7746
rect 15296 7644 15352 7654
rect 15428 7644 15489 7654
rect 15352 7588 15372 7644
rect 15428 7588 15433 7644
rect 15296 7578 15372 7588
rect 15433 7578 15489 7588
rect 15652 7644 15708 7654
rect 15708 7588 15820 7644
rect 15652 7578 15708 7588
rect 15184 7377 15260 7428
rect 14980 7084 15036 7094
rect 14980 6748 15036 7028
rect 14980 6682 15036 6692
rect 15092 6748 15148 6758
rect 14532 6570 14700 6626
rect 14868 6570 14924 6580
rect 14532 6504 14588 6514
rect 14532 6076 14588 6448
rect 14532 6010 14588 6020
rect 14644 5964 14700 6570
rect 14644 5068 14700 5908
rect 14644 5002 14700 5012
rect 14868 4956 14924 4966
rect 14980 4956 15036 4966
rect 14924 4900 14980 4956
rect 14868 4890 14924 4900
rect 14308 4778 14364 4788
rect 14308 4172 14364 4284
rect 14308 4106 14364 4116
rect 14868 4172 14924 4182
rect 14196 3098 14252 3108
rect 14420 4060 14476 4070
rect 14084 2380 14140 2996
rect 14420 2492 14476 4004
rect 14756 3948 14812 3958
rect 14756 3296 14812 3892
rect 14756 3230 14812 3240
rect 14644 3164 14700 3174
rect 14644 3052 14700 3108
rect 14644 2502 14700 2996
rect 14756 3159 14812 3169
rect 14756 3052 14812 3103
rect 14868 3052 14924 4116
rect 14812 2996 14924 3052
rect 14980 4172 15036 4900
rect 14756 2986 14812 2996
rect 14420 2426 14476 2436
rect 14532 2446 14700 2502
rect 14196 2380 14252 2390
rect 14084 2324 14196 2380
rect 14196 2314 14252 2324
rect 14532 2380 14588 2446
rect 14532 2314 14588 2324
rect 14644 2380 14700 2390
rect 14858 2380 14914 2492
rect 14980 2380 15036 4116
rect 15092 4060 15148 6692
rect 15204 5974 15260 7377
rect 15204 5908 15260 5918
rect 15316 5361 15372 7578
rect 15876 7532 15932 7680
rect 15876 7466 15932 7476
rect 15988 7420 16044 7700
rect 16100 8296 16156 8306
rect 16100 7644 16156 8240
rect 16212 7980 16268 8372
rect 16324 8362 16380 8372
rect 17220 8362 17276 8372
rect 16408 8092 16460 8148
rect 16516 8092 16616 8148
rect 16672 8092 16772 8148
rect 16828 8092 16928 8148
rect 16984 8092 17084 8148
rect 17140 8092 17192 8148
rect 16212 7914 16268 7924
rect 17332 7868 17388 7878
rect 16212 7756 16268 7766
rect 16548 7756 16604 7766
rect 16268 7700 16380 7756
rect 16212 7690 16268 7700
rect 16100 7578 16156 7588
rect 15988 7354 16044 7364
rect 15769 6987 15825 6997
rect 15647 6972 15708 6982
rect 15647 6906 15708 6916
rect 15428 6860 15484 6870
rect 15652 6819 15708 6906
rect 15764 6931 15769 6987
rect 15764 6916 15825 6931
rect 15428 5974 15484 6804
rect 15540 6748 15596 6758
rect 15540 6524 15596 6692
rect 15540 6458 15596 6468
rect 15652 6748 15708 6758
rect 15428 5918 15596 5974
rect 15428 5852 15484 5862
rect 15428 5628 15484 5796
rect 15428 5562 15484 5572
rect 15311 5296 15372 5361
rect 15428 5496 15484 5506
rect 15311 4956 15367 5296
rect 15428 5234 15484 5440
rect 15311 4697 15367 4900
rect 15423 5170 15484 5234
rect 15423 4865 15479 5170
rect 15540 5088 15596 5918
rect 15535 5078 15596 5088
rect 15591 5022 15596 5078
rect 15535 5017 15596 5022
rect 15652 5096 15708 6692
rect 15764 6748 15820 6916
rect 16212 6875 16268 6987
rect 16212 6809 16268 6819
rect 16324 6753 16380 7700
rect 16212 6697 16324 6753
rect 15764 6682 15820 6692
rect 16324 6687 16380 6697
rect 15988 6636 16044 6646
rect 15988 6514 16044 6580
rect 15988 6448 16044 6458
rect 16212 6626 16268 6636
rect 16548 6631 16604 7700
rect 16100 5964 16156 6076
rect 16100 5898 16156 5908
rect 15876 5740 15932 5852
rect 15876 5674 15932 5684
rect 16212 5628 16268 6570
rect 16324 6514 16380 6631
rect 16548 6565 16604 6575
rect 16660 6636 16716 6646
rect 16660 6524 16716 6580
rect 16660 6458 16716 6468
rect 16324 6448 16380 6458
rect 16408 6300 16460 6356
rect 16516 6300 16616 6356
rect 16672 6300 16772 6356
rect 16828 6300 16928 6356
rect 16984 6300 17084 6356
rect 17140 6300 17192 6356
rect 16660 6188 16716 6198
rect 16660 6076 16716 6132
rect 16660 6010 16716 6020
rect 16212 5562 16268 5572
rect 15652 5086 15728 5096
rect 17220 5068 17276 5078
rect 15652 5020 15728 5030
rect 15535 5012 15591 5017
rect 15652 5012 15708 5020
rect 17108 5012 17220 5068
rect 17220 5002 17276 5012
rect 15764 4956 15820 4966
rect 15540 4946 15596 4956
rect 15652 4900 15764 4956
rect 15764 4890 15820 4900
rect 15423 4808 15484 4865
rect 15311 4630 15372 4697
rect 15092 3994 15148 4004
rect 15204 4060 15260 4070
rect 14848 2324 14858 2380
rect 14914 2324 14924 2380
rect 14420 2268 14476 2278
rect 14420 2100 14476 2212
rect 14644 2268 14700 2324
rect 14766 2212 14776 2268
rect 14832 2212 14842 2268
rect 14644 2202 14700 2212
rect 14532 2156 14588 2166
rect 13972 1596 14028 1652
rect 13972 1530 14028 1540
rect 14532 1596 14588 2100
rect 14776 1959 14832 2212
rect 14532 1530 14588 1540
rect 14756 1892 14832 1959
rect 14756 1596 14812 1892
rect 14756 1530 14812 1540
rect 13402 1433 13412 1489
rect 13468 1433 13478 1489
rect 12180 746 12236 756
rect 12292 1372 12348 1382
rect 12292 1260 12348 1316
rect 12292 700 12348 1204
rect 12628 1372 12684 1382
rect 12628 1260 12684 1316
rect 12628 1194 12684 1204
rect 12740 1372 12796 1382
rect 12740 812 12796 1316
rect 12740 746 12796 756
rect 13076 1372 13132 1382
rect 12292 634 12348 644
rect 11508 522 11564 532
rect 12852 588 12908 598
rect 12908 532 13020 588
rect 12852 522 12908 532
rect 7588 476 7644 486
rect 7476 420 7588 476
rect 7364 410 7420 420
rect 7588 410 7644 420
rect 13076 476 13132 1316
rect 13412 1367 13468 1377
rect 13412 700 13468 1311
rect 13748 1372 13804 1382
rect 13412 588 13468 644
rect 13412 522 13468 532
rect 13524 588 13580 700
rect 13524 522 13580 532
rect 13748 588 13804 1316
rect 14532 1372 14588 1382
rect 14532 1204 14588 1316
rect 14980 1372 15036 2324
rect 14980 812 15036 1316
rect 15092 3276 15148 3286
rect 15092 1372 15148 3220
rect 15204 3164 15260 4004
rect 15316 3388 15372 4630
rect 15428 4396 15484 4808
rect 15428 4330 15484 4340
rect 15316 3322 15372 3332
rect 15540 3836 15596 4890
rect 16408 4508 16460 4564
rect 16516 4508 16616 4564
rect 16672 4508 16772 4564
rect 16828 4508 16928 4564
rect 16984 4508 17084 4564
rect 17140 4508 17192 4564
rect 16996 4284 17052 4294
rect 16996 4172 17052 4228
rect 16996 4106 17052 4116
rect 15316 3164 15372 3174
rect 15204 3108 15316 3164
rect 15316 3098 15372 3108
rect 15316 2380 15372 2390
rect 15204 2324 15316 2380
rect 15540 2351 15596 3780
rect 17220 3948 17276 3958
rect 17220 3836 17276 3892
rect 17220 3770 17276 3780
rect 16212 3500 16268 3510
rect 15988 3388 16044 3398
rect 15988 3220 16044 3332
rect 15652 3164 15708 3174
rect 15652 2604 15708 3108
rect 16100 3164 16156 3276
rect 16100 3098 16156 3108
rect 15652 2538 15708 2548
rect 16212 2604 16268 3444
rect 17220 3388 17276 3398
rect 17108 3332 17220 3388
rect 17220 3322 17276 3332
rect 16996 3276 17052 3286
rect 16996 3164 17052 3220
rect 16996 3098 17052 3108
rect 16408 2716 16460 2772
rect 16516 2716 16616 2772
rect 16672 2716 16772 2772
rect 16828 2716 16928 2772
rect 16984 2716 17084 2772
rect 17140 2716 17192 2772
rect 15988 2390 16044 2492
rect 15856 2380 15932 2390
rect 15316 2314 15372 2324
rect 15535 2291 15596 2351
rect 15764 2324 15856 2380
rect 15856 2314 15932 2324
rect 15988 2380 16049 2390
rect 15988 2314 16049 2324
rect 16212 2380 16268 2548
rect 16772 2604 16828 2614
rect 16212 2314 16268 2324
rect 16324 2492 16380 2502
rect 15204 2156 15260 2166
rect 15204 1708 15260 2100
rect 15535 1825 15591 2291
rect 15652 2156 15708 2166
rect 15652 2054 15708 2100
rect 15647 2044 15708 2054
rect 15784 2044 15840 2054
rect 15703 1988 15708 2044
rect 15764 1988 15784 2044
rect 15647 1978 15703 1988
rect 15764 1978 15840 1988
rect 15535 1770 15596 1825
rect 15204 1642 15260 1652
rect 15316 1484 15372 1596
rect 15316 1418 15372 1428
rect 15092 924 15148 1316
rect 15092 858 15148 868
rect 15204 1260 15260 1270
rect 14980 746 15036 756
rect 13748 522 13804 532
rect 14084 700 14140 710
rect 14084 588 14140 644
rect 15092 700 15148 710
rect 14084 522 14140 532
rect 14532 588 14588 598
rect 13076 410 13132 420
rect 14532 476 14588 532
rect 15092 588 15148 644
rect 15092 522 15148 532
rect 15204 588 15260 1204
rect 15540 1260 15596 1770
rect 15540 1194 15596 1204
rect 15204 420 15260 532
rect 15540 924 15596 934
rect 15540 476 15596 868
rect 15764 812 15820 1978
rect 15988 1367 16044 1484
rect 16212 1479 16268 1489
rect 16100 1423 16212 1479
rect 16212 1413 16268 1423
rect 16324 1479 16380 2436
rect 16324 1413 16380 1423
rect 16436 2380 16492 2390
rect 16436 1479 16492 2324
rect 16548 2380 16604 2492
rect 16548 2314 16604 2324
rect 16772 2380 16828 2548
rect 16772 2314 16828 2324
rect 17108 2604 17164 2614
rect 16772 2044 16828 2054
rect 16772 1708 16828 1988
rect 16772 1642 16828 1652
rect 17108 1596 17164 2548
rect 17108 1530 17164 1540
rect 16436 1413 16492 1423
rect 15988 1301 16044 1311
rect 16408 924 16460 980
rect 16516 924 16616 980
rect 16672 924 16772 980
rect 16828 924 16928 980
rect 16984 924 17084 980
rect 17140 924 17192 980
rect 15764 746 15820 756
rect 15876 812 15932 822
rect 14532 410 14588 420
rect 15540 410 15596 420
rect 15876 476 15932 756
rect 17332 700 17388 7812
rect 17668 7868 17724 8512
rect 17668 7802 17724 7812
rect 17892 8540 17948 8550
rect 17780 7756 17836 7766
rect 17444 7644 17500 7654
rect 17500 7588 17612 7644
rect 17444 7578 17500 7588
rect 17444 7420 17500 7430
rect 17444 6987 17500 7364
rect 17444 6916 17500 6931
rect 17780 7420 17836 7700
rect 17780 6992 17836 7364
rect 17780 6926 17836 6936
rect 17892 6870 17948 8484
rect 18228 8540 18284 8550
rect 18228 7980 18284 8484
rect 18340 8540 18396 8550
rect 18340 8372 18396 8484
rect 18676 8540 18732 9044
rect 18788 9100 18844 9380
rect 18788 9034 18844 9044
rect 19236 8876 19292 8886
rect 18676 8474 18732 8484
rect 19012 8764 19068 8774
rect 18228 7914 18284 7924
rect 18900 8316 18956 8326
rect 18228 7756 18284 7766
rect 18004 7644 18060 7654
rect 18060 7588 18172 7644
rect 18004 7578 18060 7588
rect 18004 7420 18060 7430
rect 18004 7308 18060 7364
rect 18004 7242 18060 7252
rect 17780 6814 17948 6870
rect 18004 6870 18060 6982
rect 17668 6748 17724 6758
rect 17556 6524 17612 6534
rect 17556 5964 17612 6468
rect 17556 5898 17612 5908
rect 17556 5628 17612 5638
rect 17556 4956 17612 5572
rect 17668 5516 17724 6692
rect 17668 5450 17724 5460
rect 17780 5180 17836 6814
rect 18004 6804 18060 6814
rect 17780 5114 17836 5124
rect 17892 6748 17948 6758
rect 17892 6524 17948 6692
rect 17444 4172 17500 4284
rect 17444 4106 17500 4116
rect 17444 4035 17500 4045
rect 17444 3276 17500 3979
rect 17444 3210 17500 3220
rect 17556 2380 17612 4900
rect 17892 4284 17948 6468
rect 17892 4218 17948 4228
rect 18004 5740 18060 5750
rect 17892 4060 17948 4070
rect 17780 3836 17836 3846
rect 17780 3612 17836 3780
rect 17780 3546 17836 3556
rect 17780 3276 17836 3286
rect 17780 2604 17836 3220
rect 17892 3164 17948 4004
rect 17892 3098 17948 3108
rect 18004 2736 18060 5684
rect 18116 5705 18172 7588
rect 18228 6972 18284 7700
rect 18340 7756 18396 7868
rect 18340 7690 18396 7700
rect 18676 7532 18732 7542
rect 18228 6906 18284 6916
rect 18340 7420 18396 7430
rect 18228 6636 18284 6646
rect 18228 6076 18284 6580
rect 18228 6010 18284 6020
rect 18340 5852 18396 7364
rect 18564 6636 18620 6646
rect 18564 6076 18620 6580
rect 18564 6010 18620 6020
rect 18228 5796 18340 5852
rect 18340 5786 18396 5796
rect 18116 5649 18396 5705
rect 18116 4956 18172 4966
rect 18116 4788 18172 4900
rect 18340 4172 18396 5649
rect 18564 5516 18620 5526
rect 18228 3836 18284 3846
rect 18116 3164 18172 3174
rect 18116 3032 18172 3108
rect 18228 3164 18284 3780
rect 18340 3500 18396 4116
rect 18340 3434 18396 3444
rect 18452 4732 18508 4742
rect 18228 3098 18284 3108
rect 18116 2976 18284 3032
rect 17780 2538 17836 2548
rect 17892 2680 18060 2736
rect 17556 2314 17612 2324
rect 17668 2268 17724 2278
rect 17668 2156 17724 2212
rect 17668 2090 17724 2100
rect 17556 1708 17612 1820
rect 17892 1708 17948 2680
rect 18004 2604 18060 2614
rect 18004 2492 18060 2548
rect 18228 2604 18284 2976
rect 18452 2716 18508 4676
rect 18564 3948 18620 5460
rect 18676 5068 18732 7476
rect 18900 5852 18956 8260
rect 19012 6880 19068 8708
rect 19236 8764 19292 8820
rect 19236 8698 19292 8708
rect 19124 8428 19180 8540
rect 19124 7868 19180 8372
rect 19124 7802 19180 7812
rect 19348 7644 19404 10164
rect 19796 10220 19852 10332
rect 19796 10154 19852 10164
rect 19572 9996 19628 10006
rect 19572 8764 19628 9940
rect 19684 9660 19740 9670
rect 19684 9548 19740 9604
rect 19684 9482 19740 9492
rect 20244 9314 20300 11284
rect 20580 11004 20636 11014
rect 20468 10444 20524 10454
rect 20356 10388 20468 10444
rect 20468 10378 20524 10388
rect 20244 9248 20300 9258
rect 19572 8698 19628 8708
rect 19684 9212 19740 9222
rect 19684 8540 19740 9156
rect 19684 8474 19740 8484
rect 20132 9202 20188 9212
rect 20132 8764 20188 9146
rect 19684 7868 19740 7878
rect 19684 7756 19740 7812
rect 19684 7690 19740 7700
rect 19908 7756 19964 7766
rect 19348 7420 19404 7588
rect 19908 7644 19964 7700
rect 19908 7578 19964 7588
rect 19348 7354 19404 7364
rect 19572 7532 19628 7542
rect 19012 6814 19068 6824
rect 19124 6865 19180 6977
rect 19124 6799 19180 6809
rect 18900 5786 18956 5796
rect 19012 6748 19068 6758
rect 19348 6748 19404 6758
rect 18676 5002 18732 5012
rect 18900 5715 18956 5725
rect 18788 4732 18844 4742
rect 18788 4172 18844 4676
rect 18788 4106 18844 4116
rect 18900 4060 18956 5659
rect 19012 5068 19068 6692
rect 19236 6636 19292 6748
rect 19236 6570 19292 6580
rect 19348 6524 19404 6692
rect 19460 6636 19516 6748
rect 19460 6570 19516 6580
rect 19348 6458 19404 6468
rect 19348 6300 19404 6310
rect 19012 5002 19068 5012
rect 19236 5964 19292 5974
rect 19236 4956 19292 5908
rect 19348 5964 19404 6244
rect 19348 5898 19404 5908
rect 19572 5964 19628 7476
rect 19572 5898 19628 5908
rect 19684 6748 19740 6758
rect 19684 6636 19740 6692
rect 19684 5628 19740 6580
rect 19908 6748 19964 6758
rect 19908 6188 19964 6692
rect 19908 6122 19964 6132
rect 20020 6524 20076 6534
rect 19684 5562 19740 5572
rect 20020 5068 20076 6468
rect 20020 5002 20076 5012
rect 20132 5180 20188 8708
rect 20580 8652 20636 10948
rect 20468 7092 20524 7102
rect 20351 6972 20407 6982
rect 20407 6916 20412 6972
rect 20351 6906 20412 6916
rect 20356 6748 20412 6906
rect 20356 6193 20412 6692
rect 20468 6748 20524 7036
rect 20468 6682 20524 6692
rect 20580 6636 20636 8596
rect 20692 10332 20748 12068
rect 21140 11340 21196 13972
rect 21812 13580 21868 15535
rect 22484 15596 22540 15606
rect 22372 14924 22428 14934
rect 22260 14868 22372 14924
rect 22372 14858 22428 14868
rect 22260 13916 22316 13926
rect 22148 13860 22260 13916
rect 22148 13804 22204 13860
rect 22260 13850 22316 13860
rect 22148 13738 22204 13748
rect 21812 13514 21868 13524
rect 22484 13356 22540 15540
rect 22708 15596 22764 16436
rect 22708 15530 22764 15540
rect 22932 16044 22988 16054
rect 22932 15041 22988 15988
rect 23156 15708 23212 15718
rect 23044 15652 23156 15708
rect 23044 15596 23100 15652
rect 23156 15642 23212 15652
rect 23044 15530 23100 15540
rect 22922 14985 22932 15041
rect 22988 14985 22998 15041
rect 22932 14919 22988 14929
rect 22820 14028 22876 14038
rect 22708 13972 22820 14028
rect 22820 13962 22876 13972
rect 22484 13290 22540 13300
rect 22596 13804 22652 13814
rect 22596 13224 22652 13748
rect 22932 13804 22988 14863
rect 22932 13738 22988 13748
rect 22484 13168 22652 13224
rect 21359 13132 21420 13142
rect 21496 13132 21552 13142
rect 22148 13132 22204 13142
rect 21359 13066 21420 13076
rect 21252 12012 21308 12022
rect 21252 11452 21308 11956
rect 21252 11386 21308 11396
rect 20804 11228 20860 11238
rect 20804 11004 20860 11172
rect 20804 10938 20860 10948
rect 21028 11116 21084 11126
rect 20692 8316 20748 10276
rect 20804 10444 20860 10454
rect 20804 9436 20860 10388
rect 21028 10108 21084 11060
rect 21028 10042 21084 10052
rect 21140 10332 21196 11284
rect 21364 11340 21420 13066
rect 21476 13076 21496 13132
rect 22036 13076 22148 13132
rect 21476 13066 21552 13076
rect 22148 13066 22204 13076
rect 21476 13025 21532 13066
rect 21476 12959 21532 12969
rect 21598 13020 21654 13030
rect 21476 12888 21532 12898
rect 21598 12868 21654 12964
rect 21476 12012 21532 12832
rect 21476 11946 21532 11956
rect 21588 12817 21654 12868
rect 21364 11274 21420 11284
rect 21588 11340 21644 12817
rect 21140 9660 21196 10276
rect 21140 9594 21196 9604
rect 21028 9436 21084 9446
rect 20916 9380 21028 9436
rect 20804 9202 20860 9380
rect 21028 9370 21084 9380
rect 20804 9136 20860 9146
rect 20916 9309 20972 9319
rect 20692 8250 20748 8260
rect 20916 8540 20972 9253
rect 21588 8988 21644 11284
rect 21700 12124 21756 12134
rect 21924 12124 21980 12134
rect 21812 12068 21924 12124
rect 21700 9996 21756 12068
rect 21924 12058 21980 12068
rect 22148 11457 22204 11467
rect 22036 11401 22148 11457
rect 22148 11391 22204 11401
rect 22138 11279 22148 11335
rect 22204 11279 22214 11335
rect 21700 9930 21756 9940
rect 21588 8922 21644 8932
rect 22148 8652 22204 11279
rect 22372 10444 22428 10454
rect 22372 10276 22428 10388
rect 22484 9772 22540 13168
rect 22932 13132 22988 13142
rect 22596 12908 22652 12918
rect 22596 12256 22652 12852
rect 22932 12460 22988 13076
rect 23268 12908 23324 12918
rect 23268 12684 23324 12852
rect 23268 12618 23324 12628
rect 22932 12394 22988 12404
rect 22596 12190 22652 12200
rect 22596 12119 22652 12129
rect 22596 11004 22652 12063
rect 22820 12012 22876 12022
rect 22820 11844 22876 11956
rect 22820 11228 22876 11238
rect 22708 11172 22820 11228
rect 22820 11162 22876 11172
rect 22596 10938 22652 10948
rect 23268 11116 23324 11126
rect 22596 10444 22652 10454
rect 22596 10220 22652 10388
rect 22596 10154 22652 10164
rect 22484 9706 22540 9716
rect 22260 9548 22316 9558
rect 22932 9548 22988 9660
rect 22316 9492 22428 9548
rect 22260 9482 22316 9492
rect 22148 8586 22204 8596
rect 20916 7756 20972 8484
rect 22372 8428 22428 9492
rect 22932 9482 22988 9492
rect 23268 9548 23324 11060
rect 23268 9482 23324 9492
rect 22372 8362 22428 8372
rect 23044 8540 23100 8550
rect 21476 8316 21532 8326
rect 21140 7868 21196 7980
rect 21476 7888 21532 8260
rect 21140 7802 21196 7812
rect 21364 7832 21532 7888
rect 22148 7868 22204 7878
rect 20916 7644 20972 7700
rect 20916 7578 20972 7588
rect 21364 7756 21420 7832
rect 20804 7532 20860 7542
rect 20580 6570 20636 6580
rect 20692 6748 20748 6758
rect 20692 6524 20748 6692
rect 20692 6458 20748 6468
rect 20346 6137 20356 6193
rect 20412 6137 20422 6193
rect 20356 6071 20412 6081
rect 20244 6015 20356 6071
rect 20356 6005 20412 6015
rect 20580 5180 20636 5190
rect 19236 4890 19292 4900
rect 18900 3994 18956 4004
rect 19012 4172 19068 4182
rect 18564 3276 18620 3892
rect 18564 3210 18620 3220
rect 19012 3388 19068 4116
rect 19908 4060 19964 4172
rect 19908 3994 19964 4004
rect 20020 4060 20076 4070
rect 20132 4060 20188 5124
rect 20356 5068 20412 5180
rect 20356 5002 20412 5012
rect 20580 5068 20636 5124
rect 20580 5002 20636 5012
rect 20076 4004 20188 4060
rect 20020 3994 20076 4004
rect 19012 3276 19068 3332
rect 20020 3836 20076 3846
rect 19012 3210 19068 3220
rect 19348 3276 19404 3286
rect 18452 2650 18508 2660
rect 18676 3164 18732 3174
rect 18228 2538 18284 2548
rect 18676 2604 18732 3108
rect 19348 3164 19404 3220
rect 19348 3098 19404 3108
rect 20020 3164 20076 3780
rect 20244 3612 20300 3622
rect 20244 3388 20300 3556
rect 20804 3520 20860 7476
rect 21364 6972 21420 7700
rect 21476 7756 21532 7766
rect 21476 7532 21532 7700
rect 22148 7644 22204 7812
rect 22708 7756 22764 7766
rect 22596 7700 22708 7756
rect 22708 7690 22764 7700
rect 22148 7578 22204 7588
rect 21476 7466 21532 7476
rect 21812 7532 21868 7542
rect 21364 6906 21420 6916
rect 21028 6748 21084 6758
rect 21028 6636 21084 6692
rect 21028 6570 21084 6580
rect 21588 6748 21644 6758
rect 21252 6524 21308 6534
rect 21252 6300 21308 6468
rect 21252 6234 21308 6244
rect 21588 6076 21644 6692
rect 21588 6010 21644 6020
rect 20244 3322 20300 3332
rect 20692 3464 20860 3520
rect 21028 5852 21084 5862
rect 21028 4060 21084 5796
rect 21252 5852 21308 5964
rect 21252 5786 21308 5796
rect 21700 5852 21756 5862
rect 20020 3098 20076 3108
rect 18676 2538 18732 2548
rect 18788 2940 18844 2950
rect 18788 2604 18844 2884
rect 18788 2538 18844 2548
rect 20580 2940 20636 2950
rect 18004 2426 18060 2436
rect 18340 2492 18396 2502
rect 18116 2380 18172 2390
rect 18116 2044 18172 2324
rect 18340 2380 18396 2436
rect 20580 2492 20636 2884
rect 20580 2426 20636 2436
rect 18340 2314 18396 2324
rect 18452 2380 18508 2390
rect 18788 2380 18844 2390
rect 18676 2324 18788 2380
rect 18452 2268 18508 2324
rect 18788 2314 18844 2324
rect 18452 2202 18508 2212
rect 20356 2268 20412 2278
rect 18116 1978 18172 1988
rect 19124 2156 19180 2166
rect 17892 1652 18060 1708
rect 17556 1642 17612 1652
rect 17892 1484 17948 1596
rect 17892 1418 17948 1428
rect 16660 588 16716 700
rect 17332 634 17388 644
rect 17556 1260 17612 1270
rect 17556 588 17612 1204
rect 17444 532 17556 588
rect 16660 522 16716 532
rect 17556 522 17612 532
rect 17668 812 17724 822
rect 15876 410 15932 420
rect 10164 364 10220 374
rect 5992 28 6044 84
rect 6100 28 6200 84
rect 6256 28 6356 84
rect 6412 28 6512 84
rect 6568 28 6668 84
rect 6724 28 6776 84
rect 10164 -252 10220 308
rect 14756 364 14812 374
rect 14756 -252 14812 308
rect 17668 -252 17724 756
rect 18004 28 18060 1652
rect 18228 1596 18284 1606
rect 18228 1372 18284 1540
rect 18564 1484 18620 1596
rect 18564 1418 18620 1428
rect 18116 1316 18228 1372
rect 18228 1306 18284 1316
rect 18900 700 18956 710
rect 18340 588 18396 598
rect 18900 588 18956 644
rect 18396 532 18508 588
rect 18340 522 18396 532
rect 18900 522 18956 532
rect 17892 -28 18060 28
rect 18116 476 18172 486
rect 17892 -252 17948 -28
rect 18116 -252 18172 420
rect 18564 364 18620 374
rect 18340 140 18396 150
rect 18340 -252 18396 84
rect 18564 -252 18620 308
rect 19124 140 19180 2100
rect 20244 1484 20300 1494
rect 20132 1428 20244 1484
rect 20244 1418 20300 1428
rect 20356 1260 20412 2212
rect 20468 1484 20524 1494
rect 20524 1428 20636 1484
rect 20468 1418 20524 1428
rect 20356 1194 20412 1204
rect 20692 700 20748 3464
rect 20804 3388 20860 3398
rect 20804 3276 20860 3332
rect 20804 3210 20860 3220
rect 21028 2380 21084 4004
rect 21476 4956 21532 4966
rect 21476 4060 21532 4900
rect 21700 4956 21756 5796
rect 21700 4890 21756 4900
rect 21588 4060 21644 4070
rect 21476 4004 21588 4060
rect 21476 3276 21532 4004
rect 21588 3994 21644 4004
rect 21812 3393 21868 7476
rect 22932 7532 22988 7542
rect 22036 6860 22092 6870
rect 21924 6804 22036 6860
rect 22036 6794 22092 6804
rect 22820 6748 22876 6758
rect 22820 6580 22876 6692
rect 21924 6524 21980 6534
rect 21924 5852 21980 6468
rect 22484 6188 22540 6198
rect 21924 5786 21980 5796
rect 22148 6076 22204 6086
rect 22148 4172 22204 6020
rect 22148 4106 22204 4116
rect 22260 5852 22316 5862
rect 22260 5180 22316 5796
rect 22372 5852 22428 5964
rect 22372 5786 22428 5796
rect 21476 3210 21532 3220
rect 21588 3276 21644 3388
rect 21802 3337 21812 3393
rect 21868 3337 21878 3393
rect 21924 3276 21980 3286
rect 21812 3220 21924 3276
rect 21588 3210 21644 3220
rect 21924 3210 21980 3220
rect 22148 2940 22204 2950
rect 21028 2314 21084 2324
rect 21140 2380 21196 2390
rect 20692 588 20748 644
rect 20692 522 20748 532
rect 21140 1372 21196 2324
rect 21588 1372 21644 1382
rect 21476 1316 21588 1372
rect 21140 588 21196 1316
rect 21588 1306 21644 1316
rect 21140 522 21196 532
rect 19124 74 19180 84
rect 19348 364 19404 374
rect 19348 -195 19404 308
rect 19124 -251 19404 -195
rect 19124 -252 19180 -251
rect 22148 -252 22204 2884
rect 22260 2268 22316 5124
rect 22484 5068 22540 6132
rect 22932 5404 22988 7476
rect 22932 5338 22988 5348
rect 22484 3164 22540 5012
rect 22932 4956 22988 4966
rect 22932 4844 22988 4900
rect 23044 4956 23100 8484
rect 23044 4890 23100 4900
rect 23156 7776 23212 7786
rect 22932 4778 22988 4788
rect 23044 4172 23100 4182
rect 23156 4172 23212 7720
rect 23380 7781 23436 16772
rect 23492 16492 23548 20020
rect 23604 19180 23660 19190
rect 23604 16940 23660 19124
rect 23716 17388 23772 17398
rect 23716 17164 23772 17332
rect 23716 17098 23772 17108
rect 23604 16874 23660 16884
rect 23492 16426 23548 16436
rect 23716 15596 23772 15606
rect 23604 15372 23660 15382
rect 23604 15036 23660 15316
rect 23604 14970 23660 14980
rect 23716 13132 23772 15540
rect 23716 13066 23772 13076
rect 23716 12908 23772 12918
rect 23492 12460 23548 12470
rect 23492 8769 23548 12404
rect 23716 9660 23772 12852
rect 23716 9594 23772 9604
rect 23492 8703 23548 8713
rect 23380 7715 23436 7725
rect 23492 8632 23548 8642
rect 23380 7644 23436 7654
rect 23380 6636 23436 7588
rect 23380 6570 23436 6580
rect 23492 4284 23548 8576
rect 23716 6748 23772 6758
rect 23604 6692 23716 6748
rect 23716 6682 23772 6692
rect 23716 4956 23772 4966
rect 23604 4900 23716 4956
rect 23716 4890 23772 4900
rect 23492 4218 23548 4228
rect 23100 4116 23212 4172
rect 23044 4106 23100 4116
rect 22820 4060 22876 4070
rect 22708 4004 22820 4060
rect 22820 3994 22876 4004
rect 23044 3388 23100 3398
rect 23044 3220 23100 3332
rect 23380 3276 23436 3286
rect 23268 3220 23380 3276
rect 23380 3210 23436 3220
rect 22484 3098 22540 3108
rect 22596 3164 22652 3174
rect 22596 2996 22652 3108
rect 22484 2716 22540 2726
rect 22484 2268 22540 2660
rect 22316 2212 22428 2268
rect 22260 2202 22316 2212
rect 22260 1596 22316 1606
rect 22260 1484 22316 1540
rect 22260 1418 22316 1428
rect 22372 1484 22428 2212
rect 22484 2202 22540 2212
rect 22372 476 22428 1428
rect 23716 1372 23772 1382
rect 23604 1316 23716 1372
rect 23716 1306 23772 1316
rect 22372 410 22428 420
rect 22596 476 22652 588
rect 22596 410 22652 420
<< via2 >>
rect 2548 20244 2604 20300
rect 1092 20132 1148 20188
rect 2996 20244 3052 20300
rect 868 19348 924 19404
rect 84 18447 140 18503
rect 196 18004 252 18060
rect 196 17332 252 17388
rect 196 12852 252 12908
rect 196 9940 252 9996
rect 308 10052 364 10108
rect 84 9492 140 9548
rect 756 18676 812 18732
rect 644 17332 700 17388
rect 756 15652 812 15708
rect 644 15540 700 15596
rect 1316 19236 1372 19292
rect 1876 19348 1932 19404
rect 1988 19236 2044 19292
rect 1092 15993 1148 16049
rect 1092 15871 1148 15927
rect 1988 18676 2044 18732
rect 1540 17556 1596 17612
rect 1652 18228 1708 18284
rect 1540 17108 1596 17164
rect 2100 17444 2156 17500
rect 1876 17113 1932 17169
rect 1652 16996 1708 17052
rect 1876 16996 1932 17052
rect 1652 16772 1708 16828
rect 1764 16660 1820 16716
rect 1652 15876 1708 15932
rect 2100 16660 2156 16716
rect 1652 15652 1708 15708
rect 1316 15540 1372 15596
rect 868 15408 924 15464
rect 1428 14868 1484 14924
rect 1316 14756 1372 14812
rect 1540 14308 1596 14364
rect 1092 13748 1148 13804
rect 1092 12964 1148 13020
rect 532 12292 588 12348
rect 756 12292 812 12348
rect 532 11284 588 11340
rect 420 9940 476 9996
rect 1204 12740 1260 12796
rect 1316 12292 1372 12348
rect 1092 12180 1148 12236
rect 1428 13860 1484 13916
rect 1204 11396 1260 11452
rect 1316 11172 1372 11228
rect 980 10052 1036 10108
rect 868 9828 924 9884
rect 1092 9828 1148 9884
rect 644 9370 700 9426
rect 756 9243 812 9299
rect 84 4900 140 4956
rect 420 5124 476 5180
rect 308 4340 364 4396
rect 980 9248 1036 9304
rect 980 8708 1036 8764
rect 2324 16660 2380 16716
rect 2660 17658 2716 17714
rect 2660 17444 2716 17500
rect 2558 16772 2614 16828
rect 2212 16533 2268 16589
rect 2548 16645 2604 16701
rect 2884 16553 2940 16609
rect 2772 15764 2828 15820
rect 2884 16416 2940 16472
rect 2548 15652 2604 15708
rect 1988 15092 2044 15148
rect 2436 14980 2492 15036
rect 1876 14308 1932 14364
rect 3332 20244 3388 20300
rect 3780 20132 3836 20188
rect 4116 20132 4172 20188
rect 3668 20020 3724 20076
rect 4228 20000 4284 20056
rect 3892 19236 3948 19292
rect 3444 19012 3500 19068
rect 3332 18340 3388 18396
rect 3668 18340 3724 18396
rect 3108 18024 3164 18080
rect 3240 18116 3296 18172
rect 3780 18116 3836 18172
rect 3892 18452 3948 18508
rect 3108 17887 3164 17943
rect 3556 17444 3612 17500
rect 3230 17108 3286 17164
rect 3536 16772 3592 16828
rect 3108 16670 3164 16726
rect 4116 17892 4172 17948
rect 4116 17444 4172 17500
rect 4228 17556 4284 17612
rect 3668 16660 3724 16716
rect 3544 16538 3600 16594
rect 3108 15764 3164 15820
rect 2996 15652 3052 15708
rect 2884 15540 2940 15596
rect 3220 15092 3276 15148
rect 2548 14644 2604 14700
rect 1652 14084 1708 14140
rect 4452 20244 4508 20300
rect 5012 20244 5068 20300
rect 5348 20244 5404 20300
rect 6020 20244 6076 20300
rect 4676 20132 4732 20188
rect 6356 20244 6412 20300
rect 7364 20244 7420 20300
rect 4452 19460 4508 19516
rect 4452 19236 4508 19292
rect 4564 19124 4620 19180
rect 4340 16996 4396 17052
rect 4452 18900 4508 18956
rect 6244 19908 6300 19964
rect 6044 19740 6100 19796
rect 6200 19740 6256 19796
rect 6356 19740 6412 19796
rect 6512 19740 6568 19796
rect 6668 19740 6724 19796
rect 4900 19460 4956 19516
rect 4788 19256 4844 19312
rect 4788 19124 4844 19180
rect 4676 18788 4732 18844
rect 4900 18788 4956 18844
rect 3892 16772 3948 16828
rect 4228 16772 4284 16828
rect 4116 16660 4172 16716
rect 5348 19012 5404 19068
rect 7140 19012 7196 19068
rect 6468 18900 6524 18956
rect 5796 18564 5852 18620
rect 4676 18340 4732 18396
rect 4900 18340 4956 18396
rect 4900 18228 4956 18284
rect 4564 18116 4620 18172
rect 5236 18228 5292 18284
rect 5572 18228 5628 18284
rect 5236 17668 5292 17724
rect 5124 17444 5180 17500
rect 5908 18340 5964 18396
rect 6244 18452 6300 18508
rect 6356 18452 6412 18508
rect 8820 20244 8876 20300
rect 7588 18564 7644 18620
rect 7700 18452 7756 18508
rect 6132 18228 6188 18284
rect 9380 19908 9436 19964
rect 9044 19236 9100 19292
rect 8036 18452 8092 18508
rect 6044 17948 6100 18004
rect 6200 17948 6256 18004
rect 6356 17948 6412 18004
rect 6512 17948 6568 18004
rect 6668 17948 6724 18004
rect 5684 16996 5740 17052
rect 5460 16884 5516 16940
rect 4452 16660 4508 16716
rect 4564 16548 4620 16604
rect 5348 16548 5404 16604
rect 3780 14868 3836 14924
rect 4004 14980 4060 15036
rect 2660 14420 2716 14476
rect 1876 13748 1932 13804
rect 2324 13412 2380 13468
rect 1764 12964 1820 13020
rect 1876 12292 1932 12348
rect 1652 11172 1708 11228
rect 3108 14756 3164 14812
rect 3892 14196 3948 14252
rect 3332 14084 3388 14140
rect 3108 13860 3164 13916
rect 2996 13412 3052 13468
rect 2436 12964 2492 13020
rect 2212 12068 2268 12124
rect 2436 11284 2492 11340
rect 1652 10276 1708 10332
rect 2324 10276 2380 10332
rect 1876 10164 1932 10220
rect 1428 9604 1484 9660
rect 1520 9482 1540 9538
rect 1540 9482 1576 9538
rect 3444 13300 3500 13356
rect 3332 13076 3388 13132
rect 2996 12740 3052 12796
rect 3220 12068 3276 12124
rect 2996 11284 3052 11340
rect 2996 10836 3052 10892
rect 4564 15652 4620 15708
rect 4900 15540 4956 15596
rect 4788 15204 4844 15260
rect 4452 14995 4508 15051
rect 4564 14868 4620 14924
rect 4340 14084 4396 14140
rect 4564 14420 4620 14476
rect 4228 13972 4284 14028
rect 4228 13850 4284 13906
rect 4004 13076 4060 13132
rect 4116 13300 4172 13356
rect 3556 12180 3612 12236
rect 3892 12068 3948 12124
rect 4340 13636 4396 13692
rect 5348 15540 5404 15596
rect 4900 14420 4956 14476
rect 5236 15316 5292 15372
rect 4900 14196 4956 14252
rect 5908 16660 5964 16716
rect 5796 16548 5852 16604
rect 5796 16324 5852 16380
rect 7364 17556 7420 17612
rect 7588 16772 7644 16828
rect 7364 16660 7420 16716
rect 7028 16436 7084 16492
rect 6020 16324 6076 16380
rect 6044 16156 6100 16212
rect 6200 16156 6256 16212
rect 6356 16156 6412 16212
rect 6512 16156 6568 16212
rect 6668 16156 6724 16212
rect 6356 15871 6412 15927
rect 5572 15652 5628 15708
rect 5460 15316 5516 15372
rect 6132 15652 6188 15708
rect 6356 15749 6412 15805
rect 7252 15764 7308 15820
rect 7588 15876 7644 15932
rect 7812 16660 7868 16716
rect 6020 15540 6076 15596
rect 5796 15316 5852 15372
rect 6468 15632 6524 15688
rect 7344 15316 7400 15372
rect 7481 15316 7537 15372
rect 7924 15316 7980 15372
rect 6356 14868 6412 14924
rect 7252 14644 7308 14700
rect 6804 14532 6860 14588
rect 6044 14364 6100 14420
rect 6200 14364 6256 14420
rect 6356 14364 6412 14420
rect 6512 14364 6568 14420
rect 6668 14364 6724 14420
rect 5796 14196 5852 14252
rect 6132 14196 6188 14252
rect 8148 18340 8204 18396
rect 11956 20244 12012 20300
rect 10948 20132 11004 20188
rect 12740 20132 12796 20188
rect 16460 20636 16516 20692
rect 16616 20636 16672 20692
rect 16772 20636 16828 20692
rect 16928 20636 16984 20692
rect 17084 20636 17140 20692
rect 12292 19796 12348 19852
rect 12852 19908 12908 19964
rect 10276 19124 10332 19180
rect 10388 19348 10444 19404
rect 10276 18452 10332 18508
rect 9044 17332 9100 17388
rect 8372 16660 8377 16716
rect 8377 16660 8428 16716
rect 8509 16660 8545 16716
rect 8545 16660 8565 16716
rect 8932 16660 8988 16716
rect 9044 16772 9100 16828
rect 8377 16548 8433 16604
rect 8260 15652 8316 15708
rect 8484 16436 8540 16492
rect 8148 15428 8204 15484
rect 8036 14644 8092 14700
rect 8372 14756 8428 14812
rect 7476 14084 7532 14140
rect 4788 13860 4844 13916
rect 4676 13636 4732 13692
rect 4564 13300 4620 13356
rect 4452 13188 4508 13244
rect 4228 12404 4284 12460
rect 4340 12740 4396 12796
rect 4116 12068 4172 12124
rect 2864 10388 2920 10444
rect 3001 10388 3052 10444
rect 3052 10388 3057 10444
rect 2548 9716 2604 9772
rect 1657 9492 1713 9548
rect 1871 9492 1876 9548
rect 1876 9492 1927 9548
rect 2008 9492 2044 9548
rect 2044 9492 2064 9548
rect 2212 9492 2268 9548
rect 756 4340 812 4396
rect 868 6804 924 6860
rect 1876 7588 1932 7644
rect 1876 6804 1932 6860
rect 1652 6020 1708 6076
rect 1092 5236 1148 5292
rect 1428 5236 1484 5292
rect 1092 4900 1148 4956
rect 1316 4452 1372 4508
rect 420 4116 476 4172
rect 980 4116 1036 4172
rect 868 3220 924 3276
rect 1316 3220 1372 3276
rect 1540 5012 1596 5068
rect 1876 4900 1932 4956
rect 1764 4676 1820 4732
rect 2100 4788 2156 4844
rect 2660 9487 2716 9543
rect 2660 9365 2716 9421
rect 2548 8708 2604 8764
rect 3332 10276 3388 10332
rect 3332 10052 3388 10108
rect 3220 9228 3276 9284
rect 2324 8596 2380 8652
rect 2996 8596 3052 8652
rect 2436 8484 2492 8540
rect 2324 5124 2380 5180
rect 2660 7817 2716 7873
rect 2436 5012 2492 5068
rect 2660 7680 2716 7736
rect 3108 8484 3164 8540
rect 3444 9492 3500 9548
rect 3668 9828 3724 9884
rect 3780 9492 3836 9548
rect 3892 9716 3948 9772
rect 3556 8840 3612 8896
rect 3556 8703 3612 8759
rect 3444 8036 3500 8092
rect 3444 7812 3500 7868
rect 2772 5012 2828 5068
rect 2884 6132 2940 6188
rect 2660 4900 2716 4956
rect 2996 5012 3052 5068
rect 2884 4788 2940 4844
rect 3332 5236 3388 5292
rect 3220 4900 3276 4956
rect 3556 7588 3612 7644
rect 3780 9355 3836 9411
rect 3780 8820 3836 8876
rect 3892 8260 3948 8316
rect 5572 13972 5628 14028
rect 5236 13188 5292 13244
rect 5460 13636 5516 13692
rect 4676 12292 4732 12348
rect 5348 12292 5404 12348
rect 4116 11172 4172 11228
rect 4116 10388 4172 10444
rect 5236 11956 5292 12012
rect 4676 11284 4732 11340
rect 4564 11172 4620 11228
rect 4788 11167 4844 11223
rect 4788 10836 4844 10892
rect 5236 10388 5292 10444
rect 4452 10052 4508 10108
rect 4116 9604 4172 9660
rect 4452 9604 4508 9660
rect 4228 9360 4284 9416
rect 4116 8820 4172 8876
rect 4676 9268 4732 9324
rect 4004 8372 4060 8428
rect 3444 5124 3500 5180
rect 3444 4900 3500 4956
rect 3892 8036 3948 8092
rect 2212 4676 2268 4732
rect 1876 4564 1932 4620
rect 1540 4228 1596 4284
rect 1652 4116 1708 4172
rect 308 2996 364 3052
rect 644 2996 700 3052
rect 1540 3220 1596 3276
rect 1988 3892 2044 3948
rect 1876 3220 1932 3276
rect 1652 2660 1708 2716
rect 1876 2665 1932 2721
rect 1876 2543 1932 2599
rect 2324 4116 2380 4172
rect 2212 4004 2268 4060
rect 2212 3220 2268 3276
rect 2884 4340 2940 4396
rect 2772 4228 2828 4284
rect 2660 4004 2716 4060
rect 2548 3332 2604 3388
rect 3108 4004 3164 4060
rect 2548 3108 2604 3164
rect 2996 3108 3052 3164
rect 2100 2548 2156 2604
rect 1428 1540 1484 1596
rect 1764 1652 1820 1708
rect 1204 1316 1260 1372
rect 868 756 924 812
rect 1652 980 1708 1036
rect 2324 1540 2380 1596
rect 2436 1428 2492 1484
rect 3444 3220 3500 3276
rect 4340 8427 4396 8428
rect 4340 8372 4396 8427
rect 4452 8484 4508 8540
rect 4116 8260 4172 8316
rect 6244 13972 6300 14028
rect 7364 13860 7420 13916
rect 7924 14532 7980 14588
rect 8148 14084 8204 14140
rect 5796 13193 5852 13249
rect 5796 13071 5852 13127
rect 5684 12068 5740 12124
rect 7700 13636 7756 13692
rect 7812 13860 7868 13916
rect 6020 12964 6076 13020
rect 7140 12964 7196 13020
rect 6044 12572 6100 12628
rect 6200 12572 6256 12628
rect 6356 12572 6412 12628
rect 6512 12572 6568 12628
rect 6668 12572 6724 12628
rect 6916 12068 6972 12124
rect 6244 11732 6300 11788
rect 6044 10780 6100 10836
rect 6200 10780 6256 10836
rect 6356 10780 6412 10836
rect 6512 10780 6568 10836
rect 6668 10780 6724 10836
rect 6244 10388 6300 10444
rect 6020 10164 6076 10220
rect 6804 10164 6860 10220
rect 5684 9380 5740 9436
rect 6580 9380 6636 9436
rect 7588 12190 7644 12246
rect 7476 12068 7532 12124
rect 8036 12404 8092 12460
rect 7812 12078 7868 12134
rect 7700 11956 7756 12012
rect 7924 11951 7980 12007
rect 7700 11172 7756 11228
rect 7924 11172 7980 11228
rect 7252 10164 7308 10220
rect 6044 8988 6100 9044
rect 6200 8988 6256 9044
rect 6356 8988 6412 9044
rect 6512 8988 6568 9044
rect 6668 8988 6724 9044
rect 9380 17332 9436 17388
rect 9716 17332 9772 17388
rect 9940 17220 9996 17276
rect 9716 16670 9772 16726
rect 9940 16670 9996 16726
rect 9268 16548 9324 16604
rect 9492 16553 9548 16609
rect 9156 16436 9212 16492
rect 9492 16431 9548 16487
rect 9268 15764 9324 15820
rect 9716 16436 9772 16492
rect 8708 14756 8764 14812
rect 9380 14196 9436 14252
rect 9044 13860 9100 13916
rect 8820 13748 8876 13804
rect 8372 13636 8428 13692
rect 9380 13636 9436 13692
rect 9044 13188 9100 13244
rect 8820 12740 8876 12796
rect 8596 12180 8652 12236
rect 8484 11172 8540 11228
rect 9268 12852 9324 12908
rect 9268 12516 9324 12572
rect 9156 12068 9212 12124
rect 9044 11284 9100 11340
rect 8708 11172 8764 11228
rect 8932 10164 8988 10220
rect 8148 8820 8204 8876
rect 7028 8708 7084 8764
rect 5460 8596 5516 8652
rect 5460 8148 5516 8204
rect 5796 8260 5852 8316
rect 6916 8484 6972 8540
rect 5908 8148 5964 8204
rect 5124 7812 5180 7868
rect 4228 7588 4284 7644
rect 3892 6264 3948 6320
rect 4788 7700 4844 7756
rect 5791 7588 5847 7644
rect 7252 8484 7308 8540
rect 7588 8484 7644 8540
rect 7252 7812 7308 7868
rect 5928 7588 5984 7644
rect 6916 7583 6972 7639
rect 4676 7476 4732 7532
rect 6044 7196 6100 7252
rect 6200 7196 6256 7252
rect 6356 7196 6412 7252
rect 6512 7196 6568 7252
rect 6668 7196 6724 7252
rect 5124 6804 5180 6860
rect 4676 6692 4732 6748
rect 5236 6692 5292 6748
rect 4412 6142 4468 6198
rect 3892 5592 3948 5648
rect 4004 5908 4060 5964
rect 3780 4564 3836 4620
rect 3892 5455 3948 5511
rect 4004 5012 4060 5068
rect 3668 4228 3724 4284
rect 3892 4116 3948 4172
rect 4004 4452 4060 4508
rect 3780 3892 3836 3948
rect 3556 2772 3612 2828
rect 3892 2884 3948 2940
rect 2772 1316 2828 1372
rect 3668 1652 3724 1708
rect 3556 1540 3612 1596
rect 3668 1316 3724 1372
rect 4900 6244 4956 6300
rect 5460 6244 5516 6300
rect 4544 6050 4600 6106
rect 4798 6132 4854 6188
rect 4681 6020 4737 6076
rect 4452 5796 4508 5852
rect 4452 5640 4508 5696
rect 4228 4340 4284 4396
rect 4340 5236 4396 5292
rect 4116 4208 4172 4264
rect 4564 5012 4620 5068
rect 4676 5796 4732 5852
rect 5007 5908 5012 5964
rect 5012 5908 5063 5964
rect 4788 5645 4844 5701
rect 4900 5796 4956 5852
rect 4788 5328 4844 5384
rect 4676 4890 4732 4946
rect 4564 4116 4620 4172
rect 4452 4004 4508 4060
rect 4116 3332 4172 3388
rect 4228 2996 4284 3052
rect 4228 2772 4284 2828
rect 4452 2719 4508 2775
rect 6020 6580 6076 6636
rect 6132 6468 6188 6524
rect 6916 6468 6972 6524
rect 5684 6020 5740 6076
rect 5572 5796 5628 5852
rect 5012 5236 5068 5292
rect 6044 5404 6100 5460
rect 6200 5404 6256 5460
rect 6356 5404 6412 5460
rect 6512 5404 6568 5460
rect 6668 5404 6724 5460
rect 6132 5236 6188 5292
rect 5572 5124 5628 5180
rect 5460 4900 5516 4956
rect 5684 5012 5740 5068
rect 5684 4900 5740 4956
rect 4900 4452 4956 4508
rect 5012 4778 5068 4834
rect 4900 4228 4956 4284
rect 5124 4666 5180 4722
rect 5012 3108 5068 3164
rect 4788 2884 4844 2940
rect 4676 2719 4732 2775
rect 4228 2100 4284 2156
rect 4004 1428 4060 1484
rect 4340 1316 4396 1372
rect 3108 868 3164 924
rect 6356 4900 6412 4956
rect 6244 4788 6300 4844
rect 5908 4676 5964 4732
rect 6916 4228 6972 4284
rect 5236 4116 5292 4172
rect 5684 4116 5740 4172
rect 5236 3332 5292 3388
rect 5460 2996 5516 3052
rect 5572 2324 5628 2380
rect 5012 2212 5068 2268
rect 4676 2100 4732 2156
rect 4900 1428 4956 1484
rect 4676 644 4732 700
rect 3892 532 3948 588
rect 5348 2100 5404 2156
rect 6044 3612 6100 3668
rect 6200 3612 6256 3668
rect 6356 3612 6412 3668
rect 6512 3612 6568 3668
rect 6668 3612 6724 3668
rect 5796 3332 5852 3388
rect 6244 2212 6300 2268
rect 6044 1820 6100 1876
rect 6200 1820 6256 1876
rect 6356 1820 6412 1876
rect 6512 1820 6568 1876
rect 6668 1820 6724 1876
rect 6020 1428 6076 1484
rect 6356 1316 6412 1372
rect 7364 7812 7420 7868
rect 7364 7471 7420 7527
rect 8036 8484 8092 8540
rect 7588 7700 7608 7756
rect 7608 7700 7644 7756
rect 9156 11172 9212 11228
rect 9828 15764 9884 15820
rect 10276 16548 10332 16604
rect 10052 15204 10108 15260
rect 12404 19236 12460 19292
rect 11620 19124 11676 19180
rect 11844 19124 11900 19180
rect 11060 18676 11116 18732
rect 12628 19236 12684 19292
rect 12740 19348 12796 19404
rect 10948 18340 11004 18396
rect 10836 17332 10892 17388
rect 11284 17556 11340 17612
rect 12740 17892 12796 17948
rect 12292 17556 12348 17612
rect 11620 16324 11676 16380
rect 12068 16324 12124 16380
rect 10724 15652 10780 15708
rect 11732 15652 11788 15708
rect 11508 15540 11564 15596
rect 9940 14868 9996 14924
rect 11956 15540 12012 15596
rect 11844 14888 11900 14944
rect 9492 12404 9548 12460
rect 9604 12292 9660 12348
rect 10500 14532 10556 14588
rect 10836 14532 10892 14588
rect 10052 13748 10108 13804
rect 10612 13860 10668 13916
rect 10388 13748 10444 13804
rect 10612 13188 10668 13244
rect 9828 12740 9884 12796
rect 9716 12068 9772 12124
rect 10500 12852 10556 12908
rect 10052 12292 10108 12348
rect 9604 11844 9660 11900
rect 9268 8601 9324 8657
rect 9492 8596 9548 8652
rect 9044 8484 9100 8540
rect 9156 8372 9212 8428
rect 8596 7812 8652 7868
rect 7745 7700 7801 7756
rect 8036 7700 8092 7756
rect 7700 6804 7756 6860
rect 7476 6269 7532 6325
rect 7476 6132 7532 6188
rect 7364 6015 7420 6071
rect 7588 5236 7644 5292
rect 7812 5236 7868 5292
rect 9044 7700 9100 7756
rect 9380 8484 9436 8540
rect 9716 10500 9772 10556
rect 9828 8708 9884 8764
rect 9940 10052 9996 10108
rect 8036 5129 8092 5185
rect 8372 6264 8428 6320
rect 8036 5007 8092 5063
rect 7812 4900 7868 4956
rect 7252 4788 7308 4844
rect 7364 4116 7420 4172
rect 7364 3220 7420 3276
rect 7588 4004 7644 4060
rect 7476 3108 7532 3164
rect 8596 5796 8652 5852
rect 8596 5236 8652 5292
rect 8372 4900 8428 4956
rect 8484 4676 8540 4732
rect 8484 3780 8540 3836
rect 9380 6804 9436 6860
rect 9492 6692 9548 6748
rect 9156 5684 9212 5740
rect 9156 5358 9212 5414
rect 8932 5236 8988 5292
rect 8260 3444 8316 3500
rect 8036 3332 8092 3388
rect 7924 3108 7980 3164
rect 8820 4116 8876 4172
rect 8708 3342 8764 3398
rect 8820 3780 8876 3836
rect 8708 3108 8764 3164
rect 7476 2971 7532 3027
rect 7140 1316 7196 1372
rect 7364 2436 7420 2492
rect 7700 2441 7756 2497
rect 5684 644 5740 700
rect 4900 532 4956 588
rect 1876 420 1932 476
rect 7700 2319 7756 2375
rect 7588 2197 7644 2253
rect 8036 2202 8092 2258
rect 8260 2217 8316 2273
rect 7700 1540 7756 1596
rect 8148 1316 8204 1372
rect 8484 1540 8540 1596
rect 8596 2324 8652 2380
rect 8708 2436 8764 2492
rect 8820 2324 8876 2380
rect 9716 5241 9772 5297
rect 9604 4992 9660 5048
rect 9716 5104 9772 5160
rect 8932 3220 8988 3276
rect 9268 2212 9324 2268
rect 10052 9380 10108 9436
rect 10164 11284 10220 11340
rect 10164 10276 10220 10332
rect 9940 4340 9996 4396
rect 11732 13972 11788 14028
rect 11844 14751 11900 14807
rect 12404 15652 12460 15708
rect 12516 15988 12572 16044
rect 12068 13188 12124 13244
rect 11172 12964 11228 13020
rect 11620 13076 11676 13132
rect 12180 12964 12236 13020
rect 10836 12740 10892 12796
rect 11956 12404 12012 12460
rect 10724 12180 10780 12236
rect 10612 9940 10668 9996
rect 10724 11732 10780 11788
rect 11508 12180 11564 12236
rect 11956 11732 12012 11788
rect 11284 11172 11340 11228
rect 11060 10276 11116 10332
rect 10948 9380 11004 9436
rect 10724 9156 10780 9212
rect 11732 11172 11788 11228
rect 11508 11060 11564 11116
rect 11620 10388 11676 10444
rect 11732 10500 11788 10556
rect 12404 10388 12460 10444
rect 11732 10276 11788 10332
rect 11956 10276 12012 10332
rect 11844 10144 11900 10200
rect 12180 9492 12236 9548
rect 11508 9380 11564 9436
rect 11060 8596 11116 8652
rect 11284 8708 11340 8764
rect 11956 8708 12012 8764
rect 10612 7700 10668 7756
rect 10164 7588 10220 7644
rect 11732 7140 11788 7196
rect 10612 6804 10668 6860
rect 10164 6692 10220 6748
rect 10500 6692 10556 6748
rect 10836 6580 10892 6636
rect 11732 6804 11788 6860
rect 10164 5684 10220 5740
rect 11284 5684 11340 5740
rect 10836 5012 10892 5068
rect 11396 5236 11452 5292
rect 10047 4004 10103 4060
rect 10836 4340 10892 4396
rect 10052 3337 10108 3393
rect 10276 3332 10332 3388
rect 10052 3215 10108 3271
rect 10388 2996 10444 3052
rect 9940 2324 9996 2380
rect 9604 2100 9660 2156
rect 10164 2100 10220 2156
rect 12964 17780 13020 17836
rect 13636 20020 13692 20076
rect 13300 19908 13356 19964
rect 13300 17332 13356 17388
rect 13076 17220 13132 17276
rect 13524 16772 13580 16828
rect 12852 16548 12908 16604
rect 12964 14868 13020 14924
rect 13188 14756 13244 14812
rect 12740 13972 12796 14028
rect 12740 13076 12796 13132
rect 12628 12852 12684 12908
rect 12740 12740 12796 12796
rect 12628 11172 12684 11228
rect 13300 13972 13356 14028
rect 14308 20244 14364 20300
rect 16772 20244 16828 20300
rect 14084 18676 14140 18732
rect 14868 20132 14924 20188
rect 14532 18452 14588 18508
rect 14308 18116 14364 18172
rect 14308 17220 14364 17276
rect 13636 13524 13692 13580
rect 12852 12180 12908 12236
rect 13860 15092 13916 15148
rect 16996 19348 17052 19404
rect 15652 19236 15708 19292
rect 15092 18452 15148 18508
rect 14756 18228 14812 18284
rect 14756 17444 14812 17500
rect 14420 16772 14476 16828
rect 14644 16772 14700 16828
rect 14644 14868 14700 14924
rect 14532 14089 14588 14145
rect 14084 13972 14140 14028
rect 14644 12964 14700 13020
rect 13748 12740 13804 12796
rect 13524 12404 13580 12460
rect 14980 12852 15036 12908
rect 15092 17892 15148 17948
rect 16996 19236 17052 19292
rect 17444 19236 17500 19292
rect 16772 19124 16828 19180
rect 17332 19124 17388 19180
rect 16460 18844 16516 18900
rect 16616 18844 16672 18900
rect 16772 18844 16828 18900
rect 16928 18844 16984 18900
rect 17084 18844 17140 18900
rect 16548 18676 16604 18732
rect 15428 17444 15484 17500
rect 16100 17220 16156 17276
rect 15540 16660 15596 16716
rect 15652 16548 15708 16604
rect 15316 12964 15372 13020
rect 15540 12964 15596 13020
rect 15092 12516 15148 12572
rect 15316 12516 15372 12572
rect 14868 12404 14924 12460
rect 13412 12292 13468 12348
rect 14084 12180 14140 12236
rect 15092 12180 15148 12236
rect 12964 11956 13020 12012
rect 13860 12068 13916 12124
rect 12852 11284 12908 11340
rect 13412 11172 13468 11228
rect 13524 11060 13580 11116
rect 12740 10948 12796 11004
rect 13748 10836 13804 10892
rect 12964 9492 13020 9548
rect 12740 9156 12796 9212
rect 13188 9156 13244 9212
rect 13076 7588 13132 7644
rect 12516 7028 12572 7084
rect 12740 7140 12796 7196
rect 12964 7140 13020 7196
rect 11956 6809 12012 6865
rect 12852 7028 12908 7084
rect 12516 6814 12572 6870
rect 11956 6687 12012 6743
rect 12180 5801 12236 5857
rect 11956 4788 12012 4844
rect 11508 3108 11564 3164
rect 12516 5913 12572 5969
rect 12740 5801 12796 5857
rect 12404 5572 12460 5628
rect 12740 5572 12796 5628
rect 12404 4340 12460 4396
rect 12740 4116 12796 4172
rect 13636 10388 13692 10444
rect 13748 9492 13804 9548
rect 13412 9156 13468 9212
rect 13636 9380 13692 9436
rect 14420 12068 14476 12124
rect 14756 12068 14812 12124
rect 14532 11956 14588 12012
rect 14196 11172 14252 11228
rect 14420 10948 14476 11004
rect 14308 10831 14364 10887
rect 14196 10500 14252 10556
rect 14084 10052 14140 10108
rect 14868 10388 14924 10444
rect 15092 10276 15148 10332
rect 14196 9380 14252 9436
rect 14420 9492 14476 9548
rect 13300 7700 13356 7756
rect 13412 7924 13468 7980
rect 13188 7028 13244 7084
rect 13300 6804 13356 6860
rect 12964 5913 13020 5969
rect 12964 5572 13020 5628
rect 13300 5796 13356 5852
rect 12964 4900 13020 4956
rect 12516 3220 12572 3276
rect 13636 6804 13692 6860
rect 13860 6916 13916 6972
rect 14084 7252 14140 7308
rect 14196 8820 14252 8876
rect 14532 9248 14588 9304
rect 14980 9492 15036 9548
rect 14644 8932 14700 8988
rect 14868 9360 14924 9416
rect 14756 8484 14812 8540
rect 14644 8372 14700 8428
rect 14756 7924 14812 7980
rect 14308 6580 14364 6636
rect 13636 5908 13692 5964
rect 13524 5022 13580 5078
rect 13412 4905 13468 4961
rect 13636 4900 13692 4956
rect 13300 4340 13356 4396
rect 13412 4768 13468 4824
rect 13860 4228 13916 4284
rect 12832 3108 12888 3164
rect 12969 3108 13020 3164
rect 13020 3108 13025 3164
rect 13188 3108 13244 3164
rect 12292 2884 12348 2940
rect 12964 2884 13020 2940
rect 12180 2548 12236 2604
rect 11732 2324 11788 2380
rect 10500 2212 10556 2268
rect 10388 1988 10444 2044
rect 9940 1540 9996 1596
rect 8596 1428 8652 1484
rect 9828 1316 9884 1372
rect 11060 2212 11116 2268
rect 10612 2100 10668 2156
rect 11172 1988 11228 2044
rect 12068 2212 12124 2268
rect 10500 1545 10556 1601
rect 8708 1204 8764 1260
rect 8260 980 8316 1036
rect 8708 868 8764 924
rect 9268 644 9324 700
rect 10388 644 10444 700
rect 10500 1408 10556 1464
rect 11396 532 11452 588
rect 11508 756 11564 812
rect 12292 2324 12348 2380
rect 13300 2436 13356 2492
rect 13636 1988 13692 2044
rect 13524 1540 13580 1596
rect 14756 7140 14812 7196
rect 14756 6804 14812 6860
rect 14644 6692 14700 6748
rect 15204 9626 15260 9682
rect 15540 12068 15596 12124
rect 16884 17444 16940 17500
rect 18788 20020 18844 20076
rect 20468 20244 20524 20300
rect 21140 20244 21196 20300
rect 19684 19796 19740 19852
rect 18116 19124 18172 19180
rect 18452 19348 18508 19404
rect 17444 18452 17500 18508
rect 17561 18452 17617 18508
rect 17332 17444 17388 17500
rect 16548 17220 16604 17276
rect 16460 17052 16516 17108
rect 16616 17052 16672 17108
rect 16772 17052 16828 17108
rect 16928 17052 16984 17108
rect 17084 17052 17140 17108
rect 16884 16884 16940 16940
rect 16660 16660 16716 16716
rect 15652 11844 15708 11900
rect 15764 13860 15820 13916
rect 15988 13880 16044 13936
rect 15652 11172 15708 11228
rect 15428 10500 15484 10556
rect 15428 9502 15484 9558
rect 15540 9502 15596 9558
rect 15652 9626 15708 9682
rect 15316 9156 15372 9212
rect 15092 9044 15148 9100
rect 15316 9044 15372 9100
rect 15540 9044 15596 9100
rect 15428 8932 15484 8988
rect 15988 13743 16044 13799
rect 15876 12068 15932 12124
rect 15764 8820 15820 8876
rect 17220 15540 17276 15596
rect 16460 15260 16516 15316
rect 16616 15260 16672 15316
rect 16772 15260 16828 15316
rect 16928 15260 16984 15316
rect 17084 15260 17140 15316
rect 17220 14868 17276 14924
rect 16212 14532 16268 14588
rect 16996 14532 17052 14588
rect 16436 14308 16492 14364
rect 16548 13860 16604 13916
rect 16436 13748 16492 13804
rect 19124 19348 19180 19404
rect 18788 19236 18844 19292
rect 19460 19236 19516 19292
rect 17332 13748 17388 13804
rect 17556 13748 17612 13804
rect 16460 13468 16516 13524
rect 16616 13468 16672 13524
rect 16772 13468 16828 13524
rect 16928 13468 16984 13524
rect 17084 13468 17140 13524
rect 16884 12964 16940 13020
rect 16100 11956 16156 12012
rect 16460 11676 16516 11732
rect 16616 11676 16672 11732
rect 16772 11676 16828 11732
rect 16928 11676 16984 11732
rect 17084 11676 17140 11732
rect 17108 11284 17164 11340
rect 16212 11172 16268 11228
rect 15652 8596 15708 8652
rect 14980 8260 15036 8316
rect 14980 7588 15036 7644
rect 15764 8484 15820 8540
rect 15652 8352 15708 8408
rect 16212 10948 16268 11004
rect 19012 18340 19068 18396
rect 18788 17332 18844 17388
rect 19572 17444 19628 17500
rect 18676 16889 18732 16945
rect 18676 16767 18732 16823
rect 17668 16660 17724 16716
rect 17556 13300 17612 13356
rect 17332 10948 17388 11004
rect 17444 13076 17500 13132
rect 17556 12964 17612 13020
rect 17556 12088 17612 12144
rect 17556 11951 17612 12007
rect 17556 10836 17612 10892
rect 15988 10276 16044 10332
rect 15988 9604 16044 9660
rect 16460 9884 16516 9940
rect 16616 9884 16672 9940
rect 16772 9884 16828 9940
rect 16928 9884 16984 9940
rect 17084 9884 17140 9940
rect 16212 9380 16268 9436
rect 17108 9492 17164 9548
rect 16100 8932 16156 8988
rect 16772 8932 16828 8988
rect 16324 8820 16380 8876
rect 16100 8708 16156 8764
rect 15876 7817 15932 7873
rect 17780 15988 17836 16044
rect 18340 15988 18396 16044
rect 18340 13972 18396 14028
rect 18004 12852 18060 12908
rect 18004 12292 18060 12348
rect 18564 12964 18620 13020
rect 18228 12740 18284 12796
rect 18116 12068 18172 12124
rect 18228 11172 18284 11228
rect 17668 9940 17724 9996
rect 18228 9716 18284 9772
rect 17668 9380 17724 9436
rect 18564 10948 18620 11004
rect 18788 16548 18844 16604
rect 18900 15764 18956 15820
rect 18788 14868 18844 14924
rect 18788 13748 18844 13804
rect 19012 14308 19068 14364
rect 19124 13748 19180 13804
rect 18900 11172 18956 11228
rect 19124 12964 19180 13020
rect 19460 16548 19516 16604
rect 19572 13860 19628 13916
rect 19460 13300 19516 13356
rect 19796 18116 19852 18172
rect 20356 18676 20412 18732
rect 20468 18340 20524 18396
rect 20244 17444 20300 17500
rect 20356 16660 20412 16716
rect 20468 15993 20524 16049
rect 20468 15856 20524 15912
rect 20244 15540 20300 15596
rect 19908 14980 19964 15036
rect 19908 13972 19964 14028
rect 19684 12964 19740 13020
rect 19572 12740 19628 12796
rect 20244 13076 20300 13132
rect 20132 12745 20188 12801
rect 19348 12628 19404 12684
rect 20132 12623 20188 12679
rect 19236 12068 19292 12124
rect 20244 12068 20300 12124
rect 20580 15744 20636 15800
rect 20804 19124 20860 19180
rect 21140 18452 21196 18508
rect 21364 18452 21420 18508
rect 20692 14420 20748 14476
rect 21812 19124 21868 19180
rect 21700 18564 21756 18620
rect 21476 17780 21532 17836
rect 22820 19689 22876 19745
rect 22708 19124 22764 19180
rect 22484 18452 22540 18508
rect 22932 18228 22988 18284
rect 22260 18004 22316 18060
rect 22148 17556 22204 17612
rect 21812 16772 21868 16828
rect 22036 16212 22092 16268
rect 21140 15876 21196 15932
rect 21140 14868 21196 14924
rect 20916 14644 20972 14700
rect 20804 14196 20860 14252
rect 21140 13972 21196 14028
rect 20804 13300 20860 13356
rect 20804 12964 20860 13020
rect 21028 12964 21084 13020
rect 20692 12857 20748 12913
rect 20692 12735 20748 12791
rect 20468 11956 20524 12012
rect 19908 10836 19964 10892
rect 19348 10296 19404 10352
rect 19460 10408 19516 10464
rect 19124 10164 19180 10220
rect 19348 10164 19404 10220
rect 18452 9604 18508 9660
rect 18340 9268 18396 9324
rect 17332 9044 17388 9100
rect 17658 8932 17714 8988
rect 18676 9044 18732 9100
rect 17775 8820 17831 8876
rect 17912 8820 17968 8876
rect 18136 8820 18192 8876
rect 15988 8484 16044 8540
rect 17108 8484 17164 8540
rect 16324 8372 16380 8428
rect 17220 8372 17276 8428
rect 15296 7588 15352 7644
rect 15433 7588 15489 7644
rect 15652 7588 15708 7644
rect 14980 7028 15036 7084
rect 14868 6580 14924 6636
rect 14532 6448 14588 6504
rect 14980 4900 15036 4956
rect 14308 4116 14364 4172
rect 14196 3108 14252 3164
rect 14084 2996 14140 3052
rect 14756 3240 14812 3296
rect 14644 3108 14700 3164
rect 14756 2996 14812 3052
rect 14980 4116 15036 4172
rect 14420 2436 14476 2492
rect 14532 2324 14588 2380
rect 15204 5918 15260 5974
rect 15876 7476 15932 7532
rect 16100 8240 16156 8296
rect 16460 8092 16516 8148
rect 16616 8092 16672 8148
rect 16772 8092 16828 8148
rect 16928 8092 16984 8148
rect 17084 8092 17140 8148
rect 17332 7812 17388 7868
rect 15988 7364 16044 7420
rect 15647 6916 15652 6972
rect 15652 6916 15703 6972
rect 15428 6804 15484 6860
rect 15769 6931 15825 6987
rect 15540 6468 15596 6524
rect 15652 6692 15708 6748
rect 15428 5572 15484 5628
rect 15428 5440 15484 5496
rect 15535 5022 15591 5078
rect 16212 6819 16268 6875
rect 16324 6697 16380 6753
rect 15988 6458 16044 6514
rect 16212 6570 16268 6626
rect 16100 5908 16156 5964
rect 15876 5684 15932 5740
rect 16548 6575 16604 6631
rect 16324 6458 16380 6514
rect 16660 6468 16716 6524
rect 16460 6300 16516 6356
rect 16616 6300 16672 6356
rect 16772 6300 16828 6356
rect 16928 6300 16984 6356
rect 17084 6300 17140 6356
rect 16660 6132 16716 6188
rect 16212 5572 16268 5628
rect 15672 5030 15708 5086
rect 15708 5030 15728 5086
rect 17220 5012 17276 5068
rect 15764 4900 15820 4956
rect 15092 4004 15148 4060
rect 14858 2324 14914 2380
rect 14420 2212 14476 2268
rect 14644 2212 14700 2268
rect 14776 2212 14832 2268
rect 14532 2100 14588 2156
rect 13972 1652 14028 1708
rect 14756 1540 14812 1596
rect 13412 1433 13468 1489
rect 12292 1204 12348 1260
rect 12628 1316 12684 1372
rect 12740 756 12796 812
rect 12292 644 12348 700
rect 12852 532 12908 588
rect 7588 420 7644 476
rect 13412 644 13468 700
rect 13524 532 13580 588
rect 14532 1316 14588 1372
rect 16460 4508 16516 4564
rect 16616 4508 16672 4564
rect 16772 4508 16828 4564
rect 16928 4508 16984 4564
rect 17084 4508 17140 4564
rect 16996 4228 17052 4284
rect 15540 3780 15596 3836
rect 15316 3108 15372 3164
rect 15316 2324 15372 2380
rect 17220 3780 17276 3836
rect 16212 3444 16268 3500
rect 15988 3332 16044 3388
rect 16100 3108 16156 3164
rect 17220 3332 17276 3388
rect 16996 3220 17052 3276
rect 16460 2716 16516 2772
rect 16616 2716 16672 2772
rect 16772 2716 16828 2772
rect 16928 2716 16984 2772
rect 17084 2716 17140 2772
rect 16212 2548 16268 2604
rect 15856 2324 15876 2380
rect 15876 2324 15912 2380
rect 15993 2324 16044 2380
rect 16044 2324 16049 2380
rect 16772 2548 16828 2604
rect 16324 2436 16380 2492
rect 15647 1988 15703 2044
rect 15784 1988 15840 2044
rect 15204 1652 15260 1708
rect 15316 1428 15372 1484
rect 15092 868 15148 924
rect 15204 1204 15260 1260
rect 14980 756 15036 812
rect 13748 532 13804 588
rect 14084 644 14140 700
rect 15092 644 15148 700
rect 14532 532 14588 588
rect 15540 1204 15596 1260
rect 15204 532 15260 588
rect 15540 868 15596 924
rect 16212 1423 16268 1479
rect 16548 2324 16604 2380
rect 17108 2548 17164 2604
rect 16772 1652 16828 1708
rect 16436 1423 16492 1479
rect 15988 1311 16044 1367
rect 16460 924 16516 980
rect 16616 924 16672 980
rect 16772 924 16828 980
rect 16928 924 16984 980
rect 17084 924 17140 980
rect 15876 756 15932 812
rect 17892 8484 17948 8540
rect 17780 7700 17836 7756
rect 17444 7588 17500 7644
rect 17444 6931 17500 6987
rect 17780 7364 17836 7420
rect 18340 8484 18396 8540
rect 18788 9044 18844 9100
rect 19236 8820 19292 8876
rect 19012 8708 19068 8764
rect 18228 7924 18284 7980
rect 18004 7588 18060 7644
rect 18004 7252 18060 7308
rect 18004 6814 18060 6870
rect 17556 6468 17612 6524
rect 17556 5572 17612 5628
rect 17668 5460 17724 5516
rect 17892 6468 17948 6524
rect 17444 4116 17500 4172
rect 17444 3979 17500 4035
rect 17780 3556 17836 3612
rect 17892 3108 17948 3164
rect 18340 7700 18396 7756
rect 18228 6916 18284 6972
rect 18340 7364 18396 7420
rect 18228 6020 18284 6076
rect 18564 6580 18620 6636
rect 18340 5796 18396 5852
rect 18116 4900 18172 4956
rect 18564 5460 18620 5516
rect 18228 3780 18284 3836
rect 18340 3444 18396 3500
rect 17780 2548 17836 2604
rect 17556 2324 17612 2380
rect 17668 2100 17724 2156
rect 17556 1652 17612 1708
rect 18004 2548 18060 2604
rect 19124 8372 19180 8428
rect 19796 10164 19852 10220
rect 19572 9940 19628 9996
rect 19684 9604 19740 9660
rect 20580 10948 20636 11004
rect 20468 10388 20524 10444
rect 20244 9258 20300 9314
rect 19684 9156 19740 9212
rect 20132 9146 20188 9202
rect 19684 7700 19740 7756
rect 19908 7588 19964 7644
rect 19348 7364 19404 7420
rect 19124 6809 19180 6865
rect 18900 5796 18956 5852
rect 19012 6692 19068 6748
rect 19236 6580 19292 6636
rect 19460 6580 19516 6636
rect 19348 6468 19404 6524
rect 19348 6244 19404 6300
rect 19572 5908 19628 5964
rect 19684 6580 19740 6636
rect 19908 6132 19964 6188
rect 19684 5572 19740 5628
rect 20020 5012 20076 5068
rect 20468 7036 20524 7092
rect 20351 6916 20407 6972
rect 22372 14868 22428 14924
rect 21812 13524 21868 13580
rect 22708 15540 22764 15596
rect 22932 15988 22988 16044
rect 22820 13972 22876 14028
rect 22484 13300 22540 13356
rect 22596 13748 22652 13804
rect 21359 13076 21364 13132
rect 21364 13076 21415 13132
rect 21252 11956 21308 12012
rect 21140 11284 21196 11340
rect 20804 10948 20860 11004
rect 20692 10276 20748 10332
rect 20804 10388 20860 10444
rect 21028 10052 21084 10108
rect 21496 13076 21552 13132
rect 22148 13076 22204 13132
rect 21598 12964 21654 13020
rect 21476 12832 21532 12888
rect 21364 11284 21420 11340
rect 21140 9604 21196 9660
rect 21028 9380 21084 9436
rect 20804 9146 20860 9202
rect 20916 9253 20972 9309
rect 21924 12068 21980 12124
rect 22148 11401 22204 11457
rect 22148 11279 22204 11335
rect 21700 9940 21756 9996
rect 21588 8932 21644 8988
rect 22372 10388 22428 10444
rect 23268 12628 23324 12684
rect 22596 12200 22652 12256
rect 22820 11956 22876 12012
rect 22820 11172 22876 11228
rect 22596 10948 22652 11004
rect 22596 10164 22652 10220
rect 22148 8596 22204 8652
rect 22932 9492 22988 9548
rect 23268 9492 23324 9548
rect 21140 7812 21196 7868
rect 20916 7700 20972 7756
rect 20804 7476 20860 7532
rect 20580 6580 20636 6636
rect 20692 6468 20748 6524
rect 20356 6137 20412 6193
rect 20356 6015 20412 6071
rect 20132 5124 20188 5180
rect 19236 4900 19292 4956
rect 18900 4004 18956 4060
rect 19012 4116 19068 4172
rect 19908 4004 19964 4060
rect 20356 5012 20412 5068
rect 20580 5124 20636 5180
rect 19012 3332 19068 3388
rect 20020 3780 20076 3836
rect 19348 3220 19404 3276
rect 18452 2660 18508 2716
rect 18676 3108 18732 3164
rect 20244 3556 20300 3612
rect 22708 7700 22764 7756
rect 21476 7476 21532 7532
rect 21364 6916 21420 6972
rect 21028 6580 21084 6636
rect 21252 6244 21308 6300
rect 21588 6020 21644 6076
rect 21028 5796 21084 5852
rect 21252 5796 21308 5852
rect 21700 5796 21756 5852
rect 18788 2548 18844 2604
rect 18340 2436 18396 2492
rect 20580 2436 20636 2492
rect 18788 2324 18844 2380
rect 18452 2212 18508 2268
rect 18116 1988 18172 2044
rect 17892 1428 17948 1484
rect 17332 644 17388 700
rect 17556 1204 17612 1260
rect 16660 532 16716 588
rect 17556 532 17612 588
rect 17668 756 17724 812
rect 6044 28 6100 84
rect 6200 28 6256 84
rect 6356 28 6412 84
rect 6512 28 6568 84
rect 6668 28 6724 84
rect 18228 1540 18284 1596
rect 18564 1428 18620 1484
rect 18228 1316 18284 1372
rect 18900 644 18956 700
rect 18340 532 18396 588
rect 18340 84 18396 140
rect 20244 1428 20300 1484
rect 20468 1428 20524 1484
rect 20356 1204 20412 1260
rect 20804 3332 20860 3388
rect 21476 4900 21532 4956
rect 22036 6804 22092 6860
rect 22820 6692 22876 6748
rect 22484 6132 22540 6188
rect 21924 5796 21980 5852
rect 22148 6020 22204 6076
rect 22372 5796 22428 5852
rect 22260 5124 22316 5180
rect 21812 3337 21868 3393
rect 21588 3220 21644 3276
rect 21924 3220 21980 3276
rect 20692 532 20748 588
rect 21140 1316 21196 1372
rect 21588 1316 21644 1372
rect 19124 84 19180 140
rect 22932 5348 22988 5404
rect 23044 4900 23100 4956
rect 23156 7720 23212 7776
rect 22932 4788 22988 4844
rect 23716 17108 23772 17164
rect 23604 16884 23660 16940
rect 23492 16436 23548 16492
rect 23604 15316 23660 15372
rect 23716 13076 23772 13132
rect 23716 12852 23772 12908
rect 23492 12404 23548 12460
rect 23380 7725 23436 7781
rect 23492 8576 23548 8632
rect 23380 6580 23436 6636
rect 23716 6692 23772 6748
rect 23716 4900 23772 4956
rect 22820 4004 22876 4060
rect 23044 3332 23100 3388
rect 23380 3220 23436 3276
rect 22596 3108 22652 3164
rect 22484 2660 22540 2716
rect 22260 1540 22316 1596
rect 22372 1428 22428 1484
rect 23716 1316 23772 1372
rect 22596 420 22652 476
<< metal3 >>
rect 16408 20636 16460 20692
rect 16516 20636 16616 20692
rect 16672 20636 16772 20692
rect 16828 20636 16928 20692
rect 16984 20636 17084 20692
rect 17140 20636 17192 20692
rect 3856 20300 4366 20320
rect 2538 20244 2548 20300
rect 2604 20244 2996 20300
rect 3052 20244 3062 20300
rect 3322 20244 3332 20300
rect 3388 20264 4452 20300
rect 3388 20244 3916 20264
rect 4308 20244 4452 20264
rect 4508 20244 5012 20300
rect 5068 20244 5078 20300
rect 5338 20244 5348 20300
rect 5404 20244 6020 20300
rect 6076 20244 6086 20300
rect 6346 20244 6356 20300
rect 6412 20244 7364 20300
rect 7420 20244 7430 20300
rect 8810 20244 8820 20300
rect 8876 20244 11956 20300
rect 12012 20244 12022 20300
rect 14298 20244 14308 20300
rect 14364 20244 16772 20300
rect 16828 20244 16838 20300
rect 20458 20244 20468 20300
rect 20524 20244 21140 20300
rect 21196 20244 21206 20300
rect 1082 20132 1092 20188
rect 1148 20132 3780 20188
rect 3836 20132 3846 20188
rect 4106 20132 4116 20188
rect 4172 20132 4676 20188
rect 4732 20132 4742 20188
rect 10938 20132 10948 20188
rect 11004 20132 12740 20188
rect 12796 20132 14868 20188
rect 14924 20132 14934 20188
rect 3658 20020 3668 20076
rect 3724 20056 4284 20076
rect 3724 20020 4228 20056
rect 4218 20000 4228 20020
rect 4284 20000 4294 20056
rect 13626 20020 13636 20076
rect 13692 20020 18788 20076
rect 18844 20020 18854 20076
rect 6234 19908 6244 19964
rect 6300 19908 9380 19964
rect 9436 19908 9446 19964
rect 12842 19908 12852 19964
rect 12908 19908 13300 19964
rect 13356 19908 13366 19964
rect 12282 19796 12292 19852
rect 12348 19796 19684 19852
rect 19740 19796 19750 19852
rect 5992 19740 6044 19796
rect 6100 19740 6200 19796
rect 6256 19740 6356 19796
rect 6412 19740 6512 19796
rect 6568 19740 6668 19796
rect 6724 19740 6776 19796
rect 22810 19689 22820 19745
rect 22876 19740 22886 19745
rect 22876 19689 23716 19740
rect 22820 19684 23716 19689
rect 23772 19684 23782 19740
rect 4442 19460 4452 19516
rect 4508 19460 4900 19516
rect 4956 19460 4966 19516
rect 858 19348 868 19404
rect 924 19348 1876 19404
rect 1932 19348 1942 19404
rect 10378 19348 10388 19404
rect 10444 19348 12740 19404
rect 12796 19348 12806 19404
rect 16986 19348 16996 19404
rect 17052 19348 18452 19404
rect 18508 19348 19124 19404
rect 19180 19348 19190 19404
rect 4778 19292 4788 19312
rect 1306 19236 1316 19292
rect 1372 19236 1988 19292
rect 2044 19236 2054 19292
rect 3882 19236 3892 19292
rect 3948 19236 4452 19292
rect 4508 19236 4518 19292
rect 4676 19236 4788 19292
rect 4844 19236 4854 19312
rect 9034 19236 9044 19292
rect 9100 19236 12404 19292
rect 12460 19236 12628 19292
rect 12684 19236 15652 19292
rect 15708 19236 16996 19292
rect 17052 19236 17062 19292
rect 17434 19236 17444 19292
rect 17500 19236 18788 19292
rect 18844 19236 19460 19292
rect 19516 19236 19526 19292
rect 4554 19124 4564 19180
rect 4620 19124 4788 19180
rect 4844 19124 4854 19180
rect 10266 19124 10276 19180
rect 10332 19124 11620 19180
rect 11676 19124 11844 19180
rect 11900 19124 16772 19180
rect 16828 19124 17332 19180
rect 17388 19124 18116 19180
rect 18172 19124 18182 19180
rect 20794 19124 20804 19180
rect 20860 19124 21812 19180
rect 21868 19124 22708 19180
rect 22764 19124 22774 19180
rect 3434 19012 3444 19068
rect 3500 19012 5348 19068
rect 5404 19012 7140 19068
rect 7196 19012 7206 19068
rect 4442 18900 4452 18956
rect 4508 18900 4788 18956
rect 4844 18900 6468 18956
rect 6524 18900 6534 18956
rect 16408 18844 16460 18900
rect 16516 18844 16616 18900
rect 16672 18844 16772 18900
rect 16828 18844 16928 18900
rect 16984 18844 17084 18900
rect 17140 18844 17192 18900
rect 4666 18788 4676 18844
rect 4732 18788 4900 18844
rect 4956 18788 4966 18844
rect 6024 18732 6655 18742
rect -252 18676 756 18732
rect 812 18676 822 18732
rect 1978 18676 1988 18732
rect 2044 18686 11060 18732
rect 2044 18676 6092 18686
rect 6593 18676 11060 18686
rect 11116 18676 11126 18732
rect 14074 18676 14084 18732
rect 14140 18676 16548 18732
rect 16604 18676 16614 18732
rect 20346 18676 20356 18732
rect 20412 18676 24108 18732
rect 6152 18620 6533 18630
rect 5786 18564 5796 18620
rect 5852 18574 7588 18620
rect 5852 18564 6203 18574
rect 6477 18564 7588 18574
rect 7644 18564 7654 18620
rect 21690 18564 21700 18620
rect 21756 18564 23884 18620
rect 6244 18508 6300 18518
rect -252 18503 140 18508
rect -252 18452 84 18503
rect 74 18447 84 18452
rect 140 18447 150 18503
rect 3882 18452 3892 18508
rect 3948 18452 6244 18508
rect 6244 18441 6300 18452
rect 6356 18508 6412 18518
rect 17444 18508 17500 18518
rect 6412 18452 7700 18508
rect 7756 18452 7766 18508
rect 8026 18452 8036 18508
rect 8092 18452 10276 18508
rect 10332 18452 10342 18508
rect 14522 18452 14532 18508
rect 14588 18452 15092 18508
rect 15148 18452 17444 18508
rect 6356 18442 6412 18452
rect 17444 18442 17500 18452
rect 17561 18508 17617 18518
rect 23828 18508 23884 18564
rect 17617 18452 21140 18508
rect 21196 18452 21364 18508
rect 21420 18452 21430 18508
rect 22362 18452 22372 18508
rect 22428 18452 22484 18508
rect 22540 18452 22550 18508
rect 23828 18452 24108 18508
rect 17561 18442 17617 18452
rect 3322 18340 3332 18396
rect 3388 18340 3668 18396
rect 3724 18340 4676 18396
rect 4732 18340 4742 18396
rect 4890 18340 4900 18396
rect 4956 18340 5908 18396
rect 5964 18340 5974 18396
rect 8138 18340 8148 18396
rect 8204 18340 10948 18396
rect 11004 18340 11014 18396
rect 19002 18340 19012 18396
rect 19068 18340 20468 18396
rect 20524 18340 20534 18396
rect -252 18228 308 18284
rect 364 18228 374 18284
rect 1642 18228 1652 18284
rect 1708 18228 4900 18284
rect 4956 18228 4966 18284
rect 5226 18228 5236 18284
rect 5292 18228 5572 18284
rect 5628 18228 6132 18284
rect 6188 18228 6198 18284
rect 10938 18228 10948 18284
rect 11004 18228 14756 18284
rect 14812 18228 14822 18284
rect 22922 18228 22932 18284
rect 22988 18228 24108 18284
rect 3108 18080 3164 18172
rect 3230 18116 3240 18172
rect 3296 18116 3780 18172
rect 3836 18116 4564 18172
rect 4620 18116 4630 18172
rect 14298 18116 14308 18172
rect 14364 18116 19796 18172
rect 19852 18116 19862 18172
rect -252 18004 196 18060
rect 252 18004 262 18060
rect 3098 18004 3108 18080
rect 3164 18004 3174 18080
rect 22250 18004 22260 18060
rect 22316 18004 24108 18060
rect 5992 17948 6044 18004
rect 6100 17948 6200 18004
rect 6256 17948 6356 18004
rect 6412 17948 6512 18004
rect 6568 17948 6668 18004
rect 6724 17948 6776 18004
rect 3108 17943 4116 17948
rect 3098 17887 3108 17943
rect 3164 17892 4116 17943
rect 4172 17892 4182 17948
rect 12730 17892 12740 17948
rect 12796 17892 15092 17948
rect 15148 17892 15158 17948
rect 3164 17887 3174 17892
rect -252 17826 2910 17836
rect 3400 17826 12964 17836
rect -252 17780 12964 17826
rect 13020 17780 13030 17836
rect 21466 17780 21476 17836
rect 21532 17780 24108 17836
rect 2846 17770 3460 17780
rect 3592 17714 5236 17724
rect 2650 17658 2660 17714
rect 2716 17668 5236 17714
rect 5292 17668 5302 17724
rect 2716 17658 3650 17668
rect -252 17556 1540 17612
rect 1596 17556 1606 17612
rect 4218 17556 4228 17612
rect 4284 17556 7364 17612
rect 7420 17556 7430 17612
rect 11274 17556 11284 17612
rect 11340 17556 12292 17612
rect 12348 17556 12358 17612
rect 22138 17556 22148 17612
rect 22204 17556 24108 17612
rect 2090 17444 2100 17500
rect 2156 17444 2660 17500
rect 2716 17444 2726 17500
rect 3546 17444 3556 17500
rect 3612 17444 4116 17500
rect 4172 17444 5124 17500
rect 5180 17444 5190 17500
rect 14746 17444 14756 17500
rect 14812 17444 15428 17500
rect 15484 17444 15494 17500
rect 16874 17444 16884 17500
rect 16940 17444 17332 17500
rect 17388 17444 17398 17500
rect 19562 17444 19572 17500
rect 19628 17444 20244 17500
rect 20300 17444 20310 17500
rect 186 17332 196 17388
rect 252 17332 644 17388
rect 700 17332 710 17388
rect 9034 17332 9044 17388
rect 9100 17332 9380 17388
rect 9436 17332 9446 17388
rect 9706 17332 9716 17388
rect 9772 17332 10836 17388
rect 10892 17332 13300 17388
rect 13356 17332 18788 17388
rect 18844 17332 18854 17388
rect 23706 17332 23716 17388
rect 23772 17332 24108 17388
rect 9930 17220 9940 17276
rect 9996 17220 10164 17276
rect 10220 17220 10230 17276
rect 13066 17220 13076 17276
rect 13132 17220 14308 17276
rect 14364 17220 14374 17276
rect 16090 17220 16100 17276
rect 16156 17220 16548 17276
rect 16604 17220 16614 17276
rect 1866 17164 1876 17169
rect 1530 17108 1540 17164
rect 1596 17113 1876 17164
rect 1932 17164 1942 17169
rect 1932 17113 3230 17164
rect 1596 17108 3230 17113
rect 3286 17108 3296 17164
rect 23706 17108 23716 17164
rect 23772 17108 24108 17164
rect 16408 17052 16460 17108
rect 16516 17052 16616 17108
rect 16672 17052 16772 17108
rect 16828 17052 16928 17108
rect 16984 17052 17084 17108
rect 17140 17052 17192 17108
rect 1642 16996 1652 17052
rect 1708 16996 1876 17052
rect 1932 16996 1942 17052
rect 2538 16996 2548 17052
rect 2604 16996 4340 17052
rect 4396 16996 5684 17052
rect 5740 16996 5750 17052
rect 18666 16940 18676 16945
rect 298 16884 308 16940
rect 364 16884 5460 16940
rect 5516 16884 5526 16940
rect 16874 16884 16884 16940
rect 16940 16889 18676 16940
rect 18732 16889 18742 16945
rect 16940 16884 18732 16889
rect 23594 16884 23604 16940
rect 23660 16884 24108 16940
rect 1642 16772 1652 16828
rect 1708 16772 2558 16828
rect 2614 16772 2624 16828
rect 3525 16772 3536 16828
rect 3592 16772 3602 16828
rect 3882 16772 3892 16828
rect 3948 16772 4228 16828
rect 4284 16772 4294 16828
rect 7578 16772 7588 16828
rect 7644 16772 9044 16828
rect 9100 16772 9110 16828
rect 13514 16772 13524 16828
rect 13580 16772 14420 16828
rect 14476 16772 14644 16828
rect 14700 16772 14710 16828
rect 18676 16823 21812 16828
rect 3525 16726 3581 16772
rect 18666 16767 18676 16823
rect 18732 16772 21812 16823
rect 21868 16772 21878 16828
rect 18732 16767 18742 16772
rect 1754 16660 1764 16716
rect 1820 16660 2100 16716
rect 2156 16660 2166 16716
rect 2314 16660 2324 16716
rect 2380 16706 2527 16716
rect 2380 16701 2604 16706
rect 2380 16660 2548 16701
rect 2466 16650 2548 16660
rect 2538 16645 2548 16650
rect 2604 16645 2614 16701
rect 3098 16670 3108 16726
rect 3164 16670 3581 16726
rect 3658 16660 3668 16716
rect 3724 16660 4116 16716
rect 4172 16660 4452 16716
rect 4508 16660 4518 16716
rect 5898 16660 5908 16716
rect 5964 16660 7364 16716
rect 7420 16660 7430 16716
rect 7802 16660 7812 16716
rect 7868 16660 8372 16716
rect 8428 16660 8438 16716
rect 8499 16660 8509 16716
rect 8565 16660 8932 16716
rect 8988 16660 8998 16716
rect 9706 16670 9716 16726
rect 9772 16670 9940 16726
rect 9996 16670 10006 16726
rect 15530 16660 15540 16716
rect 15596 16660 16660 16716
rect 16716 16660 17668 16716
rect 17724 16660 17734 16716
rect 20346 16660 20356 16716
rect 20412 16660 24108 16716
rect 2202 16533 2212 16589
rect 2268 16533 2548 16589
rect 2604 16533 2614 16589
rect 2874 16553 2884 16609
rect 2940 16604 2950 16609
rect 2940 16594 3507 16604
rect 2940 16553 3544 16594
rect 2884 16548 3544 16553
rect 3448 16538 3544 16548
rect 3600 16538 3610 16594
rect 4554 16548 4564 16604
rect 4620 16548 5348 16604
rect 5404 16548 5796 16604
rect 5852 16548 5862 16604
rect 8367 16548 8377 16604
rect 8433 16548 9268 16604
rect 9324 16548 9334 16604
rect 9482 16553 9492 16609
rect 9548 16604 9558 16609
rect 9548 16553 10276 16604
rect 9492 16548 10276 16553
rect 10332 16548 10342 16604
rect 12842 16548 12852 16604
rect 12908 16548 15652 16604
rect 15708 16548 15718 16604
rect 18778 16548 18788 16604
rect 18844 16548 19460 16604
rect 19516 16548 19526 16604
rect 2884 16482 3354 16492
rect 3991 16482 7028 16492
rect 2884 16472 7028 16482
rect 2874 16416 2884 16472
rect 2940 16436 7028 16472
rect 7084 16436 8484 16492
rect 8540 16436 9156 16492
rect 9212 16487 9548 16492
rect 9212 16436 9492 16487
rect 2940 16416 2950 16436
rect 3292 16426 4048 16436
rect 9482 16431 9492 16436
rect 9548 16431 9558 16487
rect 9706 16436 9716 16492
rect 9772 16436 10948 16492
rect 11004 16436 11014 16492
rect 23482 16436 23492 16492
rect 23548 16436 24108 16492
rect 5786 16324 5796 16380
rect 5852 16324 6020 16380
rect 6076 16324 6086 16380
rect 11610 16324 11620 16380
rect 11676 16324 12068 16380
rect 12124 16324 12134 16380
rect 22026 16212 22036 16268
rect 22092 16212 24108 16268
rect 5992 16156 6044 16212
rect 6100 16156 6200 16212
rect 6256 16156 6356 16212
rect 6412 16156 6512 16212
rect 6568 16156 6668 16212
rect 6724 16156 6776 16212
rect 1082 15993 1092 16049
rect 1148 16044 1158 16049
rect 20458 16044 20468 16049
rect 1148 15993 12516 16044
rect 1092 15988 12516 15993
rect 12572 15988 17780 16044
rect 17836 15988 18340 16044
rect 18396 15993 20468 16044
rect 20524 15993 20534 16049
rect 18396 15988 20524 15993
rect 22922 15988 22932 16044
rect 22988 15988 24108 16044
rect 1092 15927 1652 15932
rect 1082 15871 1092 15927
rect 1148 15876 1652 15927
rect 1708 15876 1718 15932
rect 1148 15871 1158 15876
rect 6346 15871 6356 15927
rect 6412 15922 6422 15927
rect 6652 15922 7588 15932
rect 6412 15876 7588 15922
rect 7644 15876 7654 15932
rect 20468 15912 21140 15932
rect 6412 15871 6714 15876
rect 6356 15866 6714 15871
rect 20458 15856 20468 15912
rect 20524 15876 21140 15912
rect 21196 15876 21206 15932
rect 20524 15856 20534 15876
rect 2762 15764 2772 15820
rect 2828 15764 3108 15820
rect 3164 15764 3174 15820
rect 6778 15810 7252 15820
rect 6356 15805 7252 15810
rect 6346 15749 6356 15805
rect 6412 15764 7252 15805
rect 7308 15764 7318 15820
rect 9258 15764 9268 15820
rect 9324 15764 9828 15820
rect 9884 15764 9894 15820
rect 18890 15764 18900 15820
rect 18956 15800 20323 15820
rect 18956 15764 20580 15800
rect 6412 15754 6832 15764
rect 6412 15749 6422 15754
rect 20251 15744 20580 15764
rect 20636 15744 20646 15800
rect 23706 15764 23716 15820
rect 23772 15764 24108 15820
rect 746 15652 756 15708
rect 812 15652 1652 15708
rect 1708 15652 2548 15708
rect 2604 15652 2996 15708
rect 3052 15652 3062 15708
rect 4554 15652 4564 15708
rect 4620 15652 5572 15708
rect 5628 15652 6132 15708
rect 6188 15688 6230 15708
rect 6188 15652 6468 15688
rect 6162 15632 6468 15652
rect 6524 15632 6534 15688
rect 8250 15652 8260 15708
rect 8316 15652 10724 15708
rect 10780 15652 11732 15708
rect 11788 15652 12404 15708
rect 12460 15652 12470 15708
rect 634 15540 644 15596
rect 700 15540 1316 15596
rect 1372 15540 2884 15596
rect 2940 15540 2950 15596
rect 4890 15540 4900 15596
rect 4956 15540 5348 15596
rect 5404 15540 6020 15596
rect 6076 15540 6086 15596
rect 11498 15540 11508 15596
rect 11564 15540 11956 15596
rect 12012 15540 12022 15596
rect 17210 15540 17220 15596
rect 17276 15540 20244 15596
rect 20300 15540 20310 15596
rect 22698 15540 22708 15596
rect 22764 15540 24108 15596
rect 1130 15464 8148 15484
rect 858 15408 868 15464
rect 924 15428 8148 15464
rect 8204 15428 8214 15484
rect 924 15408 1191 15428
rect 5226 15316 5236 15372
rect 5292 15316 5460 15372
rect 5516 15316 5526 15372
rect 5786 15316 5796 15372
rect 5852 15316 7344 15372
rect 7400 15316 7410 15372
rect 7471 15316 7481 15372
rect 7537 15316 7924 15372
rect 7980 15316 7990 15372
rect 23594 15316 23604 15372
rect 23660 15316 24108 15372
rect 16408 15260 16460 15316
rect 16516 15260 16616 15316
rect 16672 15260 16772 15316
rect 16828 15260 16928 15316
rect 16984 15260 17084 15316
rect 17140 15260 17192 15316
rect 4778 15204 4788 15260
rect 4844 15204 10052 15260
rect 10108 15204 10118 15260
rect 1978 15092 1988 15148
rect 2044 15092 3220 15148
rect 3276 15092 3286 15148
rect 13850 15092 13860 15148
rect 13916 15092 21028 15148
rect 21084 15092 24108 15148
rect 4442 15036 4452 15051
rect 2426 14980 2436 15036
rect 2492 14980 4004 15036
rect 4060 14995 4452 15036
rect 4508 14995 4518 15051
rect 4060 14980 4508 14995
rect 19898 14980 19908 15036
rect 19964 14980 23884 15036
rect 11834 14924 11844 14944
rect 1418 14868 1428 14924
rect 1484 14868 3780 14924
rect 3836 14868 4564 14924
rect 4620 14868 6356 14924
rect 6412 14868 6422 14924
rect 9930 14868 9940 14924
rect 9996 14888 11844 14924
rect 11900 14888 11910 14944
rect 23828 14924 23884 14980
rect 9996 14868 11900 14888
rect 12954 14868 12964 14924
rect 13020 14868 14644 14924
rect 14700 14868 17220 14924
rect 17276 14868 18788 14924
rect 18844 14868 18854 14924
rect 21130 14868 21140 14924
rect 21196 14868 22372 14924
rect 22428 14868 22438 14924
rect 23828 14868 24108 14924
rect 1306 14756 1316 14812
rect 1372 14756 3108 14812
rect 3164 14756 3174 14812
rect 8362 14756 8372 14812
rect 8428 14756 8708 14812
rect 8764 14756 8774 14812
rect 11844 14807 13188 14812
rect 11834 14751 11844 14807
rect 11900 14756 13188 14807
rect 13244 14756 13254 14812
rect 11900 14751 11910 14756
rect 2538 14644 2548 14700
rect 2604 14644 7252 14700
rect 7308 14644 8036 14700
rect 8092 14644 8102 14700
rect 20906 14644 20916 14700
rect 20972 14644 24108 14700
rect 6794 14532 6804 14588
rect 6860 14532 7924 14588
rect 7980 14532 7990 14588
rect 10490 14532 10500 14588
rect 10556 14532 10836 14588
rect 10892 14532 10902 14588
rect 16202 14532 16212 14588
rect 16268 14532 16996 14588
rect 17052 14532 17062 14588
rect 2650 14420 2660 14476
rect 2716 14420 4564 14476
rect 4620 14420 4900 14476
rect 4956 14420 4966 14476
rect 20682 14420 20692 14476
rect 20748 14420 24108 14476
rect 5992 14364 6044 14420
rect 6100 14364 6200 14420
rect 6256 14364 6356 14420
rect 6412 14364 6512 14420
rect 6568 14364 6668 14420
rect 6724 14364 6776 14420
rect 1530 14308 1540 14364
rect 1596 14308 1876 14364
rect 1932 14308 1942 14364
rect 16426 14308 16436 14364
rect 16492 14308 19012 14364
rect 19068 14308 19078 14364
rect 3882 14196 3892 14252
rect 3948 14196 4900 14252
rect 4956 14196 4966 14252
rect 5786 14196 5796 14252
rect 5852 14196 6132 14252
rect 6188 14196 9380 14252
rect 9436 14196 9446 14252
rect 20794 14196 20804 14252
rect 20860 14196 24108 14252
rect 14522 14140 14532 14145
rect 1642 14084 1652 14140
rect 1708 14084 3332 14140
rect 3388 14084 4340 14140
rect 4396 14084 7476 14140
rect 7532 14084 8148 14140
rect 8204 14084 8214 14140
rect 14410 14084 14420 14140
rect 14476 14089 14532 14140
rect 14588 14089 14598 14145
rect 14476 14084 14588 14089
rect 3108 13916 3164 14028
rect 4218 13972 4228 14028
rect 4284 13972 5572 14028
rect 5628 13972 6244 14028
rect 6300 13972 6310 14028
rect 11722 13972 11732 14028
rect 11788 13972 12740 14028
rect 12796 13972 13300 14028
rect 13356 13972 14084 14028
rect 14140 13972 14150 14028
rect 18330 13972 18340 14028
rect 18396 13972 19908 14028
rect 19964 13972 21140 14028
rect 21196 13972 21206 14028
rect 22810 13972 22820 14028
rect 22876 13972 24108 14028
rect 15978 13916 15988 13936
rect 1418 13860 1428 13916
rect 1484 13860 3108 13916
rect 3164 13860 3174 13916
rect 4359 13911 4788 13916
rect 4228 13906 4788 13911
rect 4218 13850 4228 13906
rect 4284 13860 4788 13906
rect 4844 13860 4854 13916
rect 7354 13860 7364 13916
rect 7420 13860 7812 13916
rect 7868 13860 7878 13916
rect 9034 13860 9044 13916
rect 9100 13860 10612 13916
rect 10668 13860 10678 13916
rect 15754 13860 15764 13916
rect 15820 13880 15988 13916
rect 16044 13880 16054 13936
rect 15820 13860 16044 13880
rect 16538 13860 16548 13916
rect 16604 13860 19572 13916
rect 19628 13860 19638 13916
rect 4284 13855 4417 13860
rect 4284 13850 4294 13855
rect 1082 13748 1092 13804
rect 1148 13748 1876 13804
rect 1932 13748 1942 13804
rect 8810 13748 8820 13804
rect 8876 13748 10052 13804
rect 10108 13748 10388 13804
rect 10444 13748 10454 13804
rect 15988 13799 16436 13804
rect 15978 13743 15988 13799
rect 16044 13748 16436 13799
rect 16492 13748 16502 13804
rect 17322 13748 17332 13804
rect 17388 13748 17556 13804
rect 17612 13748 17622 13804
rect 18778 13748 18788 13804
rect 18844 13748 19124 13804
rect 19180 13748 19190 13804
rect 22586 13748 22596 13804
rect 22652 13748 24108 13804
rect 16044 13743 16054 13748
rect 4330 13636 4340 13692
rect 4396 13636 4676 13692
rect 4732 13636 5460 13692
rect 5516 13636 5526 13692
rect 7690 13636 7700 13692
rect 7756 13636 8372 13692
rect 8428 13636 9380 13692
rect 9436 13636 9446 13692
rect 13626 13524 13636 13580
rect 13692 13524 13702 13580
rect 21802 13524 21812 13580
rect 21868 13524 24108 13580
rect 2314 13412 2324 13468
rect 2380 13412 2996 13468
rect 3052 13412 4844 13468
rect 13636 13412 13692 13524
rect 16408 13468 16460 13524
rect 16516 13468 16616 13524
rect 16672 13468 16772 13524
rect 16828 13468 16928 13524
rect 16984 13468 17084 13524
rect 17140 13468 17192 13524
rect 4788 13356 4844 13412
rect 5646 13356 6000 13361
rect 3434 13300 3444 13356
rect 3500 13300 4116 13356
rect 4172 13300 4564 13356
rect 4620 13300 4630 13356
rect 4788 13305 17556 13356
rect 4788 13300 5706 13305
rect 5942 13300 17556 13305
rect 17612 13300 17622 13356
rect 19450 13300 19460 13356
rect 19516 13300 20804 13356
rect 20860 13300 20870 13356
rect 22474 13300 22484 13356
rect 22540 13300 24108 13356
rect 4442 13188 4452 13244
rect 4508 13188 5236 13244
rect 5292 13188 5302 13244
rect 5786 13193 5796 13249
rect 5852 13244 5862 13249
rect 5852 13193 9044 13244
rect 5796 13188 9044 13193
rect 9100 13188 9110 13244
rect 10602 13188 10612 13244
rect 10668 13188 12068 13244
rect 12124 13188 12134 13244
rect 3322 13076 3332 13132
rect 3388 13076 4004 13132
rect 4060 13127 5852 13132
rect 4060 13076 5796 13127
rect 5786 13071 5796 13076
rect 5852 13071 5862 13127
rect 11610 13076 11620 13132
rect 11676 13076 11732 13132
rect 11788 13076 11798 13132
rect 12730 13076 12740 13132
rect 12796 13076 17444 13132
rect 17500 13076 17510 13132
rect 20234 13076 20244 13132
rect 20300 13076 21359 13132
rect 21415 13076 21425 13132
rect 21486 13076 21496 13132
rect 21552 13076 22148 13132
rect 22204 13076 22214 13132
rect 23706 13076 23716 13132
rect 23772 13076 24108 13132
rect 1082 12964 1092 13020
rect 1148 12964 1764 13020
rect 1820 12964 2436 13020
rect 2492 12964 2502 13020
rect 6010 12964 6020 13020
rect 6076 12964 7140 13020
rect 7196 12964 7206 13020
rect 11162 12964 11172 13020
rect 11228 12964 12180 13020
rect 12236 12964 12246 13020
rect 14634 12964 14644 13020
rect 14700 12964 15316 13020
rect 15372 12964 15382 13020
rect 15530 12964 15540 13020
rect 15596 12964 16884 13020
rect 16940 12964 16950 13020
rect 17546 12964 17556 13020
rect 17612 12964 18564 13020
rect 18620 12964 18630 13020
rect 19114 12964 19124 13020
rect 19180 12964 19684 13020
rect 19740 12964 19750 13020
rect 20794 12964 20804 13020
rect 20860 12964 21028 13020
rect 21084 12964 21598 13020
rect 21654 12964 21664 13020
rect 186 12852 196 12908
rect 252 12852 9268 12908
rect 9324 12852 9334 12908
rect 10490 12852 10500 12908
rect 10556 12852 12628 12908
rect 12684 12852 12694 12908
rect 14970 12852 14980 12908
rect 15036 12852 17668 12908
rect 17724 12852 18004 12908
rect 18060 12852 18070 12908
rect 20682 12857 20692 12913
rect 20748 12908 20758 12913
rect 20748 12888 21532 12908
rect 20748 12857 21476 12888
rect 20692 12852 21476 12857
rect 21466 12832 21476 12852
rect 21532 12832 21542 12888
rect 23706 12852 23716 12908
rect 23772 12852 24108 12908
rect 20122 12796 20132 12801
rect 1194 12740 1204 12796
rect 1260 12740 1428 12796
rect 1484 12740 2996 12796
rect 3052 12740 4340 12796
rect 4396 12740 8820 12796
rect 8876 12740 8886 12796
rect 9818 12740 9828 12796
rect 9884 12740 10836 12796
rect 10892 12740 12740 12796
rect 12796 12740 13748 12796
rect 13804 12740 18228 12796
rect 18284 12740 18294 12796
rect 19562 12740 19572 12796
rect 19628 12745 20132 12796
rect 20188 12796 20198 12801
rect 20188 12791 20748 12796
rect 20188 12745 20692 12791
rect 19628 12740 20692 12745
rect 20682 12735 20692 12740
rect 20748 12735 20758 12791
rect 19338 12628 19348 12684
rect 19404 12679 20188 12684
rect 19404 12628 20132 12679
rect 5992 12572 6044 12628
rect 6100 12572 6200 12628
rect 6256 12572 6356 12628
rect 6412 12572 6512 12628
rect 6568 12572 6668 12628
rect 6724 12572 6776 12628
rect 20122 12623 20132 12628
rect 20188 12623 20198 12679
rect 23258 12628 23268 12684
rect 23324 12628 24108 12684
rect 9258 12516 9268 12572
rect 9324 12516 15092 12572
rect 15148 12516 15316 12572
rect 15372 12516 15382 12572
rect 4218 12404 4228 12460
rect 4284 12404 8036 12460
rect 8092 12404 9492 12460
rect 9548 12404 9558 12460
rect 11946 12404 11956 12460
rect 12012 12404 13524 12460
rect 13580 12404 14868 12460
rect 14924 12404 14934 12460
rect 23482 12404 23492 12460
rect 23548 12404 24108 12460
rect 522 12292 532 12348
rect 588 12292 756 12348
rect 812 12292 1316 12348
rect 1372 12292 1876 12348
rect 1932 12292 1942 12348
rect 4666 12292 4676 12348
rect 4732 12292 5348 12348
rect 5404 12292 5414 12348
rect 9594 12292 9604 12348
rect 9660 12292 10052 12348
rect 10108 12292 10118 12348
rect 13402 12292 13412 12348
rect 13468 12292 18004 12348
rect 18060 12292 18070 12348
rect 1082 12180 1092 12236
rect 1148 12180 3556 12236
rect 3612 12180 3622 12236
rect 7578 12190 7588 12246
rect 7644 12236 8325 12246
rect 7644 12190 8596 12236
rect 8264 12180 8596 12190
rect 8652 12180 8662 12236
rect 10714 12180 10724 12236
rect 10780 12180 11508 12236
rect 11564 12180 11574 12236
rect 12842 12180 12852 12236
rect 12908 12180 14084 12236
rect 14140 12180 15092 12236
rect 15148 12180 15158 12236
rect 22586 12200 22596 12256
rect 22652 12236 22662 12256
rect 22652 12200 24108 12236
rect 22596 12180 24108 12200
rect 2202 12068 2212 12124
rect 2268 12068 3220 12124
rect 3276 12068 3892 12124
rect 3948 12068 3958 12124
rect 4106 12068 4116 12124
rect 4172 12068 5684 12124
rect 5740 12068 5750 12124
rect 6906 12068 6916 12124
rect 6972 12068 7476 12124
rect 7532 12068 7542 12124
rect 7802 12078 7812 12134
rect 7868 12129 7878 12134
rect 7868 12124 8184 12129
rect 17546 12124 17556 12144
rect 7868 12078 9156 12124
rect 7812 12073 9156 12078
rect 8124 12068 9156 12073
rect 9212 12068 9716 12124
rect 9772 12068 9782 12124
rect 13850 12068 13860 12124
rect 13916 12068 14420 12124
rect 14476 12068 14486 12124
rect 14746 12068 14756 12124
rect 14812 12068 15540 12124
rect 15596 12068 15606 12124
rect 15866 12068 15876 12124
rect 15932 12088 17556 12124
rect 17612 12088 17622 12144
rect 15932 12068 17612 12088
rect 18106 12068 18116 12124
rect 18172 12068 19236 12124
rect 19292 12068 20244 12124
rect 20300 12068 21924 12124
rect 21980 12068 21990 12124
rect 5226 11956 5236 12012
rect 5292 11956 7700 12012
rect 7756 12007 7980 12012
rect 7756 11956 7924 12007
rect 7914 11951 7924 11956
rect 7980 11951 7990 12007
rect 12954 11956 12964 12012
rect 13020 11956 14532 12012
rect 14588 11956 14598 12012
rect 16090 11956 16100 12012
rect 16156 12007 17612 12012
rect 16156 11956 17556 12007
rect 17546 11951 17556 11956
rect 17612 11951 17622 12007
rect 20010 11956 20020 12012
rect 20076 11956 20468 12012
rect 20524 11956 20534 12012
rect 21242 11956 21252 12012
rect 21308 11956 22372 12012
rect 22428 11956 22820 12012
rect 22876 11956 22886 12012
rect 9594 11844 9604 11900
rect 9660 11844 15652 11900
rect 15708 11844 15718 11900
rect 6234 11732 6244 11788
rect 6300 11732 10724 11788
rect 10780 11732 11956 11788
rect 12012 11732 12022 11788
rect 16408 11676 16460 11732
rect 16516 11676 16616 11732
rect 16672 11676 16772 11732
rect 16828 11676 16928 11732
rect 16984 11676 17084 11732
rect 17140 11676 17192 11732
rect 1194 11396 1204 11452
rect 1260 11396 1428 11452
rect 1484 11396 1494 11452
rect 22138 11401 22148 11457
rect 22204 11452 22214 11457
rect 22204 11401 24108 11452
rect 22148 11396 24108 11401
rect 522 11284 532 11340
rect 588 11284 2436 11340
rect 2492 11284 2996 11340
rect 3052 11284 3062 11340
rect 4666 11284 4676 11340
rect 4732 11284 9044 11340
rect 9100 11284 9110 11340
rect 10154 11284 10164 11340
rect 10220 11284 12852 11340
rect 12908 11284 12918 11340
rect 17098 11284 17108 11340
rect 17164 11284 21140 11340
rect 21196 11284 21206 11340
rect 21354 11284 21364 11340
rect 21420 11335 22204 11340
rect 21420 11284 22148 11335
rect 22138 11279 22148 11284
rect 22204 11279 22214 11335
rect 1306 11172 1316 11228
rect 1372 11172 1652 11228
rect 1708 11172 1718 11228
rect 4106 11172 4116 11228
rect 4172 11172 4564 11228
rect 4620 11172 4630 11228
rect 4788 11223 7700 11228
rect 4778 11167 4788 11223
rect 4844 11172 7700 11223
rect 7756 11172 7924 11228
rect 7980 11172 8484 11228
rect 8540 11172 8550 11228
rect 8698 11172 8708 11228
rect 8764 11172 9156 11228
rect 9212 11172 9222 11228
rect 11274 11172 11284 11228
rect 11340 11172 11732 11228
rect 11788 11172 11798 11228
rect 12618 11172 12628 11228
rect 12684 11172 13412 11228
rect 13468 11172 14196 11228
rect 14252 11172 14262 11228
rect 15642 11172 15652 11228
rect 15708 11172 16212 11228
rect 16268 11172 16278 11228
rect 18218 11172 18228 11228
rect 18284 11172 18900 11228
rect 18956 11172 18966 11228
rect 22810 11172 22820 11228
rect 22876 11172 24108 11228
rect 4844 11167 4854 11172
rect 11498 11060 11508 11116
rect 11564 11060 13524 11116
rect 13580 11060 13590 11116
rect 12730 10948 12740 11004
rect 12796 10948 14420 11004
rect 14476 10948 14980 11004
rect 15036 10948 15046 11004
rect 16202 10948 16212 11004
rect 16268 10948 17332 11004
rect 17388 10948 17398 11004
rect 18554 10948 18564 11004
rect 18620 10948 20580 11004
rect 20636 10948 20804 11004
rect 20860 10948 22596 11004
rect 22652 10948 22662 11004
rect 2986 10836 2996 10892
rect 3052 10836 4788 10892
rect 4844 10836 4854 10892
rect 13738 10836 13748 10892
rect 13804 10887 14364 10892
rect 13804 10836 14308 10887
rect 5992 10780 6044 10836
rect 6100 10780 6200 10836
rect 6256 10780 6356 10836
rect 6412 10780 6512 10836
rect 6568 10780 6668 10836
rect 6724 10780 6776 10836
rect 14298 10831 14308 10836
rect 14364 10831 14374 10887
rect 17546 10836 17556 10892
rect 17612 10836 19908 10892
rect 19964 10836 19974 10892
rect 9706 10500 9716 10556
rect 9772 10500 11732 10556
rect 11788 10500 11798 10556
rect 14186 10500 14196 10556
rect 14252 10500 15428 10556
rect 15484 10500 15494 10556
rect 19191 10444 19460 10464
rect 2538 10388 2548 10444
rect 2604 10388 2864 10444
rect 2920 10388 2930 10444
rect 2991 10388 3001 10444
rect 3057 10388 4116 10444
rect 4172 10388 4182 10444
rect 5226 10388 5236 10444
rect 5292 10388 6244 10444
rect 6300 10388 6310 10444
rect 11610 10388 11620 10444
rect 11676 10388 12404 10444
rect 12460 10388 13636 10444
rect 13692 10388 13702 10444
rect 14858 10388 14868 10444
rect 14924 10388 18564 10444
rect 18620 10408 19460 10444
rect 19516 10444 19943 10464
rect 19516 10408 20468 10444
rect 18620 10388 19246 10408
rect 19877 10388 20468 10408
rect 20524 10388 20534 10444
rect 20794 10388 20804 10444
rect 20860 10388 22372 10444
rect 22428 10388 22438 10444
rect 1642 10276 1652 10332
rect 1708 10276 2324 10332
rect 2380 10276 3332 10332
rect 3388 10276 3398 10332
rect 10154 10276 10164 10332
rect 10220 10276 11060 10332
rect 11116 10276 11126 10332
rect 11722 10276 11732 10332
rect 11788 10276 11956 10332
rect 12012 10276 12022 10332
rect 15082 10276 15092 10332
rect 15148 10276 15988 10332
rect 16044 10276 16054 10332
rect 19338 10296 19348 10352
rect 19404 10342 19414 10352
rect 19404 10332 19778 10342
rect 19404 10296 20692 10332
rect 19348 10286 20692 10296
rect 19348 10276 19404 10286
rect 19717 10276 20692 10286
rect 20748 10276 20758 10332
rect 1866 10164 1876 10220
rect 1932 10164 6020 10220
rect 6076 10164 6804 10220
rect 6860 10164 7252 10220
rect 7308 10164 8932 10220
rect 8988 10164 8998 10220
rect 11722 10164 11732 10220
rect 11788 10200 11900 10220
rect 11788 10164 11844 10200
rect 11834 10144 11844 10164
rect 11900 10144 11910 10200
rect 19114 10164 19124 10220
rect 19180 10164 19348 10220
rect 19404 10164 19414 10220
rect 19786 10164 19796 10220
rect 19852 10164 22596 10220
rect 22652 10164 22662 10220
rect 298 10052 308 10108
rect 364 10052 980 10108
rect 1036 10052 3332 10108
rect 3388 10052 3398 10108
rect 4442 10052 4452 10108
rect 4508 10052 9940 10108
rect 9996 10052 10006 10108
rect 14074 10052 14084 10108
rect 14140 10052 21028 10108
rect 21084 10052 21094 10108
rect 186 9940 196 9996
rect 252 9940 420 9996
rect 476 9940 10612 9996
rect 10668 9940 10678 9996
rect 17658 9940 17668 9996
rect 17724 9940 19572 9996
rect 19628 9940 21700 9996
rect 21756 9940 21766 9996
rect 16408 9884 16460 9940
rect 16516 9884 16616 9940
rect 16672 9884 16772 9940
rect 16828 9884 16928 9940
rect 16984 9884 17084 9940
rect 17140 9884 17192 9940
rect 858 9828 868 9884
rect 924 9828 1092 9884
rect 1148 9828 3668 9884
rect 3724 9828 3734 9884
rect 2538 9716 2548 9772
rect 2604 9716 3892 9772
rect 3948 9716 3958 9772
rect 15194 9738 15204 9794
rect 15260 9772 16014 9794
rect 15260 9738 18228 9772
rect 15956 9718 18228 9738
rect 15957 9716 18228 9718
rect 18284 9716 18294 9772
rect 1418 9604 1428 9660
rect 1484 9604 4116 9660
rect 4172 9604 4452 9660
rect 4508 9604 4518 9660
rect 15194 9626 15204 9682
rect 15260 9626 15428 9682
rect 15484 9626 15652 9682
rect 15708 9626 15718 9682
rect 15978 9604 15988 9660
rect 16044 9604 18452 9660
rect 18508 9604 18518 9660
rect 19674 9604 19684 9660
rect 19740 9604 21140 9660
rect 21196 9604 21252 9660
rect 21308 9604 21318 9660
rect 15428 9558 15484 9570
rect 15223 9548 15428 9558
rect 74 9492 84 9548
rect 140 9538 1464 9548
rect 140 9492 1520 9538
rect 1395 9482 1520 9492
rect 1576 9482 1586 9538
rect 1647 9492 1657 9548
rect 1713 9492 1871 9548
rect 1927 9492 1937 9548
rect 1998 9492 2008 9548
rect 2064 9492 2212 9548
rect 2268 9492 2278 9548
rect 2708 9543 3444 9548
rect 2650 9487 2660 9543
rect 2716 9492 3444 9543
rect 3500 9492 3780 9548
rect 3836 9492 3846 9548
rect 12170 9492 12180 9548
rect 12236 9492 12964 9548
rect 13020 9492 13030 9548
rect 13738 9492 13748 9548
rect 13804 9492 14420 9548
rect 14476 9492 14486 9548
rect 14970 9492 14980 9548
rect 15036 9502 15428 9548
rect 15036 9492 15281 9502
rect 15428 9492 15484 9502
rect 15540 9558 15596 9568
rect 15596 9548 15810 9558
rect 15596 9502 17108 9548
rect 15540 9492 15596 9502
rect 15754 9492 17108 9502
rect 17164 9492 17174 9548
rect 22922 9492 22932 9548
rect 22988 9492 23268 9548
rect 23324 9492 23334 9548
rect 2716 9487 2824 9492
rect 2660 9482 2824 9487
rect 873 9426 1343 9436
rect 1735 9426 2442 9436
rect 634 9370 644 9426
rect 700 9421 2716 9426
rect 700 9380 2660 9421
rect 700 9370 928 9380
rect 1279 9370 1793 9380
rect 2380 9370 2660 9380
rect 2650 9365 2660 9370
rect 2716 9365 2726 9421
rect 3780 9411 4228 9416
rect 3770 9355 3780 9411
rect 3836 9360 4228 9411
rect 4284 9360 4294 9416
rect 5674 9380 5684 9436
rect 5740 9380 6580 9436
rect 6636 9380 6646 9436
rect 10042 9380 10052 9436
rect 10108 9380 10948 9436
rect 11004 9380 11014 9436
rect 11498 9380 11508 9436
rect 11564 9380 13636 9436
rect 13692 9380 13702 9436
rect 14186 9380 14196 9436
rect 14252 9416 16212 9436
rect 14252 9380 14868 9416
rect 14858 9360 14868 9380
rect 14924 9380 16212 9416
rect 16268 9380 16278 9436
rect 17658 9380 17668 9436
rect 17724 9380 21028 9436
rect 21084 9380 21094 9436
rect 14924 9360 14934 9380
rect 3836 9355 3846 9360
rect 756 9299 980 9304
rect 746 9243 756 9299
rect 812 9248 980 9299
rect 1036 9248 1046 9304
rect 4431 9284 4676 9324
rect 812 9243 822 9248
rect 3210 9228 3220 9284
rect 3276 9268 4676 9284
rect 4732 9268 4742 9324
rect 15061 9304 18340 9324
rect 3276 9228 4495 9268
rect 14522 9248 14532 9304
rect 14588 9268 18340 9304
rect 18396 9268 18406 9324
rect 14588 9248 15136 9268
rect 20234 9258 20244 9314
rect 20300 9309 20972 9314
rect 20300 9258 20916 9309
rect 20906 9253 20916 9258
rect 20972 9253 20982 9309
rect 10714 9156 10724 9212
rect 10780 9156 12740 9212
rect 12796 9156 13188 9212
rect 13244 9156 13412 9212
rect 13468 9156 13478 9212
rect 15306 9156 15316 9212
rect 15372 9156 19684 9212
rect 19740 9156 19750 9212
rect 20122 9146 20132 9202
rect 20188 9146 20804 9202
rect 20860 9146 20870 9202
rect 15082 9044 15092 9100
rect 15148 9044 15316 9100
rect 15372 9044 15382 9100
rect 15530 9044 15540 9100
rect 15596 9044 17332 9100
rect 17388 9044 18676 9100
rect 18732 9044 18788 9100
rect 18844 9044 18854 9100
rect 5992 8988 6044 9044
rect 6100 8988 6200 9044
rect 6256 8988 6356 9044
rect 6412 8988 6512 9044
rect 6568 8988 6668 9044
rect 6724 8988 6776 9044
rect 14634 8932 14644 8988
rect 14700 8932 15428 8988
rect 15484 8932 15494 8988
rect 16090 8932 16100 8988
rect 16156 8932 16772 8988
rect 16828 8932 16838 8988
rect 17648 8932 17658 8988
rect 17714 8932 21588 8988
rect 21644 8932 21654 8988
rect 3546 8840 3556 8896
rect 3612 8876 3622 8896
rect 3612 8840 3780 8876
rect 3556 8820 3780 8840
rect 3836 8820 3846 8876
rect 4106 8820 4116 8876
rect 4172 8820 8148 8876
rect 8204 8820 8214 8876
rect 14186 8820 14196 8876
rect 14252 8820 15764 8876
rect 15820 8820 15830 8876
rect 16314 8820 16324 8876
rect 16380 8820 17775 8876
rect 17831 8820 17841 8876
rect 17902 8820 17912 8876
rect 17968 8820 18060 8876
rect 18126 8820 18136 8876
rect 18192 8820 19236 8876
rect 19292 8820 19302 8876
rect 970 8708 980 8764
rect 1036 8708 2548 8764
rect 2604 8708 2614 8764
rect 3556 8759 7028 8764
rect 3546 8703 3556 8759
rect 3612 8708 7028 8759
rect 7084 8708 7094 8764
rect 9818 8708 9828 8764
rect 9884 8708 11284 8764
rect 11340 8708 11956 8764
rect 12012 8708 12022 8764
rect 16090 8708 16100 8764
rect 16156 8708 17668 8764
rect 17724 8708 19012 8764
rect 19068 8708 19078 8764
rect 3612 8703 3622 8708
rect 2314 8596 2324 8652
rect 2380 8596 2996 8652
rect 3052 8596 3062 8652
rect 4330 8596 4340 8652
rect 4396 8596 5460 8652
rect 5516 8596 5526 8652
rect 9258 8601 9268 8657
rect 9324 8652 9334 8657
rect 9324 8601 9492 8652
rect 9268 8596 9492 8601
rect 9548 8596 9558 8652
rect 11050 8596 11060 8652
rect 11116 8596 11620 8652
rect 11676 8596 11686 8652
rect 15642 8596 15652 8652
rect 15708 8596 22148 8652
rect 22204 8596 22214 8652
rect 23492 8632 23716 8652
rect 23482 8576 23492 8632
rect 23548 8596 23716 8632
rect 23772 8596 23782 8652
rect 23548 8576 23558 8596
rect 2426 8484 2436 8540
rect 2492 8484 3108 8540
rect 3164 8484 3174 8540
rect 4442 8484 4452 8540
rect 4508 8484 6916 8540
rect 6972 8484 6982 8540
rect 7242 8484 7252 8540
rect 7308 8484 7588 8540
rect 7644 8484 8036 8540
rect 8092 8484 8102 8540
rect 9034 8484 9044 8540
rect 9100 8484 9380 8540
rect 9436 8484 9446 8540
rect 14410 8484 14420 8540
rect 14476 8484 14756 8540
rect 14812 8484 14822 8540
rect 15754 8484 15764 8540
rect 15820 8484 15988 8540
rect 16044 8484 16054 8540
rect 17098 8484 17108 8540
rect 17164 8484 17892 8540
rect 17948 8484 18340 8540
rect 18396 8484 18406 8540
rect 3994 8372 4004 8428
rect 4060 8372 4340 8428
rect 4396 8372 9156 8428
rect 9212 8372 9222 8428
rect 14634 8372 14644 8428
rect 14700 8408 15708 8428
rect 14700 8372 15652 8408
rect 15642 8352 15652 8372
rect 15708 8352 15718 8408
rect 16314 8372 16324 8428
rect 16380 8372 17220 8428
rect 17276 8372 19124 8428
rect 19180 8372 19190 8428
rect 3882 8260 3892 8316
rect 3948 8260 4116 8316
rect 4172 8260 4182 8316
rect 5450 8260 5460 8316
rect 5516 8260 5796 8316
rect 5852 8260 5862 8316
rect 14970 8260 14980 8316
rect 15036 8296 15563 8316
rect 15036 8260 16100 8296
rect 15500 8240 16100 8260
rect 16156 8240 16166 8296
rect 5450 8148 5460 8204
rect 5516 8148 5908 8204
rect 5964 8148 5974 8204
rect 16408 8092 16460 8148
rect 16516 8092 16616 8148
rect 16672 8092 16772 8148
rect 16828 8092 16928 8148
rect 16984 8092 17084 8148
rect 17140 8092 17192 8148
rect 3434 8036 3444 8092
rect 3500 8036 3892 8092
rect 3948 8036 3958 8092
rect 13402 7924 13412 7980
rect 13468 7924 14756 7980
rect 14812 7924 15204 7980
rect 15260 7924 15270 7980
rect 17322 7924 17332 7980
rect 17388 7924 18228 7980
rect 18284 7924 18294 7980
rect 2650 7817 2660 7873
rect 2716 7868 2726 7873
rect 2716 7817 3444 7868
rect 2660 7812 3444 7817
rect 3500 7812 3510 7868
rect 5114 7812 5124 7868
rect 5180 7812 7252 7868
rect 7308 7812 7364 7868
rect 7420 7812 8596 7868
rect 8652 7812 8662 7868
rect 15866 7817 15876 7873
rect 15932 7868 15942 7873
rect 15932 7817 17332 7868
rect 15876 7812 17332 7817
rect 17388 7812 17398 7868
rect 21018 7812 21028 7868
rect 21084 7812 21140 7868
rect 21196 7812 21206 7868
rect 23370 7776 23380 7781
rect 2660 7736 4788 7756
rect 2650 7680 2660 7736
rect 2716 7700 4788 7736
rect 4844 7700 7588 7756
rect 7644 7700 7654 7756
rect 7735 7700 7745 7756
rect 7801 7700 8036 7756
rect 8092 7700 8102 7756
rect 9034 7700 9044 7756
rect 9100 7700 10612 7756
rect 10668 7700 10678 7756
rect 13290 7700 13300 7756
rect 13356 7700 17332 7756
rect 17388 7700 17398 7756
rect 17770 7700 17780 7756
rect 17836 7700 18340 7756
rect 18396 7700 19684 7756
rect 19740 7700 19750 7756
rect 20906 7700 20916 7756
rect 20972 7700 22708 7756
rect 22764 7700 22774 7756
rect 23146 7720 23156 7776
rect 23212 7725 23380 7776
rect 23436 7725 23446 7781
rect 23212 7720 23436 7725
rect 2716 7680 2726 7700
rect 1866 7588 1876 7644
rect 1932 7624 2539 7644
rect 2920 7624 3556 7644
rect 1932 7588 3556 7624
rect 3612 7588 3622 7644
rect 4218 7588 4228 7644
rect 4284 7588 5791 7644
rect 5847 7588 5857 7644
rect 5918 7588 5928 7644
rect 5984 7639 6972 7644
rect 5984 7588 6916 7639
rect 2474 7568 2987 7588
rect 6906 7583 6916 7588
rect 6972 7583 6982 7639
rect 10154 7588 10164 7644
rect 10220 7588 13076 7644
rect 13132 7588 13142 7644
rect 14970 7588 14980 7644
rect 15036 7588 15296 7644
rect 15352 7588 15362 7644
rect 15423 7588 15433 7644
rect 15489 7588 15652 7644
rect 15708 7588 17444 7644
rect 17500 7588 18004 7644
rect 18060 7588 19908 7644
rect 19964 7588 19974 7644
rect 4666 7476 4676 7532
rect 4732 7476 4900 7532
rect 4956 7527 6748 7532
rect 4956 7476 7364 7527
rect 6683 7471 7364 7476
rect 7420 7471 7430 7527
rect 15866 7476 15876 7532
rect 15932 7476 20804 7532
rect 20860 7476 21476 7532
rect 21532 7476 21542 7532
rect 15978 7364 15988 7420
rect 16044 7364 17780 7420
rect 17836 7364 17846 7420
rect 18330 7364 18340 7420
rect 18396 7364 19348 7420
rect 19404 7364 19414 7420
rect 14074 7252 14084 7308
rect 14140 7252 18004 7308
rect 18060 7252 18070 7308
rect 5992 7196 6044 7252
rect 6100 7196 6200 7252
rect 6256 7196 6356 7252
rect 6412 7196 6512 7252
rect 6568 7196 6668 7252
rect 6724 7196 6776 7252
rect 11722 7140 11732 7196
rect 11788 7140 12740 7196
rect 12796 7140 12806 7196
rect 12954 7140 12964 7196
rect 13020 7140 14756 7196
rect 14812 7140 14822 7196
rect 12506 7028 12516 7084
rect 12572 7028 12852 7084
rect 12908 7028 12918 7084
rect 13178 7028 13188 7084
rect 13244 7028 14980 7084
rect 15036 7028 15046 7084
rect 20458 7036 20468 7092
rect 20524 7036 20817 7092
rect 15769 6987 15825 6997
rect 13850 6916 13860 6972
rect 13916 6916 15647 6972
rect 15703 6916 15713 6972
rect 15825 6931 17444 6987
rect 17500 6931 17510 6987
rect 18749 6972 19522 6977
rect 20761 6972 20817 7036
rect 15769 6916 15825 6931
rect 18218 6916 18228 6972
rect 18284 6921 20351 6972
rect 18284 6916 18818 6921
rect 19459 6916 20351 6921
rect 20407 6916 20417 6972
rect 20761 6916 21364 6972
rect 21420 6916 21430 6972
rect 11946 6860 11956 6865
rect 858 6804 868 6860
rect 924 6804 1876 6860
rect 1932 6804 1942 6860
rect 5114 6804 5124 6860
rect 5180 6804 7700 6860
rect 7756 6804 7766 6860
rect 9370 6804 9380 6860
rect 9436 6804 10612 6860
rect 10668 6804 11732 6860
rect 11788 6809 11956 6860
rect 12012 6809 12022 6865
rect 12506 6814 12516 6870
rect 12572 6860 12693 6870
rect 12572 6814 13300 6860
rect 11788 6804 12012 6809
rect 12635 6804 13300 6814
rect 13356 6804 13636 6860
rect 13692 6804 13702 6860
rect 14746 6804 14756 6860
rect 14812 6804 14980 6860
rect 15036 6804 15046 6860
rect 15418 6804 15428 6860
rect 15484 6804 15596 6860
rect 16202 6819 16212 6875
rect 16268 6870 16278 6875
rect 16268 6819 18004 6870
rect 16212 6814 18004 6819
rect 18060 6814 18070 6870
rect 19114 6809 19124 6865
rect 19180 6860 19395 6865
rect 19180 6809 22036 6860
rect 19331 6804 22036 6809
rect 22092 6804 22102 6860
rect 15942 6748 16324 6753
rect 4666 6692 4676 6748
rect 4732 6692 5236 6748
rect 5292 6692 5302 6748
rect 9482 6692 9492 6748
rect 9548 6692 10164 6748
rect 10220 6692 10500 6748
rect 10556 6692 10566 6748
rect 11956 6743 14644 6748
rect 11946 6687 11956 6743
rect 12012 6692 14644 6743
rect 14700 6692 14710 6748
rect 15642 6692 15652 6748
rect 15708 6697 16324 6748
rect 16380 6697 16390 6753
rect 19012 6748 19278 6753
rect 15708 6692 16002 6697
rect 19002 6692 19012 6748
rect 19068 6697 20020 6748
rect 19068 6692 19078 6697
rect 19217 6692 20020 6697
rect 20076 6692 22820 6748
rect 22876 6692 22886 6748
rect 23706 6692 23716 6748
rect 23772 6692 24108 6748
rect 12012 6687 12022 6692
rect 6010 6580 6020 6636
rect 6076 6580 10836 6636
rect 10892 6580 10902 6636
rect 14298 6580 14308 6636
rect 14364 6580 14868 6636
rect 14924 6580 14934 6636
rect 16212 6626 16548 6631
rect 16202 6570 16212 6626
rect 16268 6575 16548 6626
rect 16604 6575 16614 6631
rect 18554 6580 18564 6636
rect 18620 6580 19236 6636
rect 19292 6580 19460 6636
rect 19516 6580 19526 6636
rect 19674 6580 19684 6636
rect 19740 6580 20580 6636
rect 20636 6580 21028 6636
rect 21084 6580 23380 6636
rect 23436 6580 23446 6636
rect 16268 6570 16278 6575
rect 6122 6468 6132 6524
rect 6188 6468 6916 6524
rect 6972 6468 6982 6524
rect 14978 6504 15540 6524
rect 14522 6448 14532 6504
rect 14588 6468 15540 6504
rect 15596 6468 15606 6524
rect 14588 6448 15042 6468
rect 15978 6458 15988 6514
rect 16044 6458 16324 6514
rect 16380 6458 16390 6514
rect 16650 6468 16660 6524
rect 16716 6468 17332 6524
rect 17388 6468 17556 6524
rect 17612 6468 17622 6524
rect 17882 6468 17892 6524
rect 17948 6468 19348 6524
rect 19404 6468 20692 6524
rect 20748 6468 20758 6524
rect 3882 6264 3892 6320
rect 3948 6300 4759 6320
rect 3948 6264 4900 6300
rect 4697 6244 4900 6264
rect 4956 6244 5460 6300
rect 5516 6244 5526 6300
rect 7466 6269 7476 6325
rect 7532 6320 7542 6325
rect 7532 6269 8372 6320
rect 7476 6264 8372 6269
rect 8428 6264 8438 6320
rect 16408 6300 16460 6356
rect 16516 6300 16616 6356
rect 16672 6300 16772 6356
rect 16828 6300 16928 6356
rect 16984 6300 17084 6356
rect 17140 6300 17192 6356
rect 20160 6300 20716 6305
rect 19338 6244 19348 6300
rect 19404 6249 21252 6300
rect 19404 6244 20227 6249
rect 20640 6244 21252 6249
rect 21308 6244 21318 6300
rect 4250 6188 4412 6198
rect 2874 6132 2884 6188
rect 2940 6142 4412 6188
rect 4468 6142 4478 6198
rect 7476 6188 7532 6193
rect 2940 6132 4312 6142
rect 4788 6132 4798 6188
rect 4854 6132 7476 6188
rect 7532 6132 7542 6188
rect 16650 6132 16660 6188
rect 16716 6132 19908 6188
rect 19964 6132 19974 6188
rect 20346 6137 20356 6193
rect 20412 6188 20422 6193
rect 20412 6137 22484 6188
rect 20356 6132 22484 6137
rect 22540 6132 22550 6188
rect 4534 6086 4544 6106
rect 4452 6076 4544 6086
rect 1642 6020 1652 6076
rect 1708 6050 4544 6076
rect 4600 6050 4610 6106
rect 1708 6030 4600 6050
rect 1708 6020 4518 6030
rect 4671 6020 4681 6076
rect 4737 6020 5684 6076
rect 5740 6071 9044 6076
rect 5740 6020 7364 6071
rect 7354 6015 7364 6020
rect 7420 6020 9044 6071
rect 9100 6020 9110 6076
rect 18218 6020 18228 6076
rect 18284 6071 21588 6076
rect 18284 6020 20356 6071
rect 7420 6015 7430 6020
rect 20346 6015 20356 6020
rect 20412 6020 21588 6071
rect 21644 6020 22148 6076
rect 22204 6020 22214 6076
rect 20412 6015 20422 6020
rect 3994 5908 4004 5964
rect 4060 5908 5007 5964
rect 5063 5908 5073 5964
rect 12506 5913 12516 5969
rect 12572 5913 12964 5969
rect 13020 5913 13030 5969
rect 14911 5964 15204 5974
rect 13626 5908 13636 5964
rect 13692 5918 15204 5964
rect 15260 5964 15806 5974
rect 15260 5918 16100 5964
rect 13692 5908 14970 5918
rect 15745 5908 16100 5918
rect 16156 5908 19572 5964
rect 19628 5908 19638 5964
rect 4442 5796 4452 5852
rect 4508 5796 4676 5852
rect 4732 5796 4742 5852
rect 4890 5796 4900 5852
rect 4956 5796 5572 5852
rect 5628 5796 8596 5852
rect 8652 5796 8662 5852
rect 12170 5801 12180 5857
rect 12236 5801 12740 5857
rect 12796 5801 12806 5857
rect 21252 5852 21308 5964
rect 13290 5796 13300 5852
rect 13356 5796 18004 5852
rect 18060 5847 18211 5852
rect 18330 5847 18340 5852
rect 18060 5796 18340 5847
rect 18396 5796 18406 5852
rect 18778 5796 18788 5852
rect 18844 5796 18900 5852
rect 18956 5796 18966 5852
rect 21018 5796 21028 5852
rect 21084 5796 21252 5852
rect 21308 5796 21700 5852
rect 21756 5796 21766 5852
rect 21914 5796 21924 5852
rect 21980 5796 22372 5852
rect 22428 5796 22438 5852
rect 18148 5791 18396 5796
rect 4452 5696 4508 5706
rect 4778 5696 4788 5701
rect 3882 5628 3892 5648
rect 3770 5572 3780 5628
rect 3836 5592 3892 5628
rect 3948 5592 3958 5648
rect 4508 5645 4788 5696
rect 4844 5645 4854 5701
rect 9146 5684 9156 5740
rect 9212 5684 10164 5740
rect 10220 5684 10230 5740
rect 11274 5684 11284 5740
rect 11340 5684 15876 5740
rect 15932 5684 15942 5740
rect 4508 5640 4844 5645
rect 4452 5630 4508 5640
rect 3836 5572 3948 5592
rect 12394 5572 12404 5628
rect 12460 5572 12740 5628
rect 12796 5572 12806 5628
rect 12954 5572 12964 5628
rect 13020 5572 15428 5628
rect 15484 5572 16212 5628
rect 16268 5572 17556 5628
rect 17612 5572 19684 5628
rect 19740 5572 19750 5628
rect 3892 5511 4335 5516
rect 3882 5455 3892 5511
rect 3948 5460 4335 5511
rect 4391 5460 4401 5516
rect 15674 5496 17668 5516
rect 3948 5455 3958 5460
rect 5992 5404 6044 5460
rect 6100 5404 6200 5460
rect 6256 5404 6356 5460
rect 6412 5404 6512 5460
rect 6568 5404 6668 5460
rect 6724 5404 6776 5460
rect 15418 5440 15428 5496
rect 15484 5460 17668 5496
rect 17724 5460 18564 5516
rect 18620 5460 18630 5516
rect 15484 5440 15734 5460
rect 4788 5384 5460 5404
rect 4778 5328 4788 5384
rect 4844 5348 5460 5384
rect 5516 5348 5526 5404
rect 9146 5358 9156 5414
rect 9212 5404 10388 5414
rect 9212 5358 13636 5404
rect 10328 5348 13636 5358
rect 13692 5384 15169 5404
rect 15800 5384 22932 5404
rect 13692 5348 22932 5384
rect 22988 5348 22998 5404
rect 4844 5328 4854 5348
rect 15106 5328 15860 5348
rect 7878 5292 8276 5297
rect 1082 5236 1092 5292
rect 1148 5236 1428 5292
rect 1484 5236 3332 5292
rect 3388 5236 4340 5292
rect 4396 5236 4406 5292
rect 5002 5236 5012 5292
rect 5068 5236 6132 5292
rect 6188 5236 7588 5292
rect 7644 5236 7812 5292
rect 7868 5241 8596 5292
rect 7868 5236 7934 5241
rect 8216 5236 8596 5241
rect 8652 5236 8932 5292
rect 8988 5236 8998 5292
rect 9706 5241 9716 5297
rect 9772 5292 9782 5297
rect 9772 5241 11396 5292
rect 9716 5236 11396 5241
rect 11452 5236 11462 5292
rect 410 5124 420 5180
rect 476 5124 2324 5180
rect 2380 5124 2390 5180
rect 3434 5124 3444 5180
rect 3500 5124 5572 5180
rect 5628 5124 5638 5180
rect 8026 5129 8036 5185
rect 8092 5180 8102 5185
rect 8092 5160 9772 5180
rect 8092 5129 9716 5160
rect 8036 5124 9716 5129
rect 9706 5104 9716 5124
rect 9772 5104 9782 5160
rect 15535 5078 15591 5180
rect 20122 5124 20132 5180
rect 20188 5124 20580 5180
rect 20636 5124 22260 5180
rect 22316 5124 22326 5180
rect 12967 5068 13524 5078
rect 1530 5012 1540 5068
rect 1596 5012 2436 5068
rect 2492 5012 2502 5068
rect 2762 5012 2772 5068
rect 2828 5012 2996 5068
rect 3052 5012 4004 5068
rect 4060 5012 4070 5068
rect 4472 5012 4564 5068
rect 4620 5012 4630 5068
rect 5674 5012 5684 5068
rect 5740 5063 8092 5068
rect 5740 5012 8036 5063
rect 8026 5007 8036 5012
rect 8092 5007 8102 5063
rect 9919 5048 10836 5068
rect 9594 4992 9604 5048
rect 9660 5012 10836 5048
rect 10892 5022 13524 5068
rect 13580 5022 13590 5078
rect 10892 5012 13027 5022
rect 15525 5017 15535 5078
rect 15591 5017 15601 5078
rect 15662 5030 15672 5086
rect 15728 5068 15738 5086
rect 15728 5030 17220 5068
rect 15672 5012 17220 5030
rect 17276 5012 17286 5068
rect 20010 5012 20020 5068
rect 20076 5012 20356 5068
rect 20412 5012 20422 5068
rect 9660 4992 9983 5012
rect 13402 4956 13412 4961
rect 74 4900 84 4956
rect 140 4900 1092 4956
rect 1148 4900 1158 4956
rect 1866 4900 1876 4956
rect 1932 4900 2660 4956
rect 2716 4900 2726 4956
rect 3210 4900 3220 4956
rect 3276 4900 3444 4956
rect 3500 4900 3510 4956
rect 4778 4951 4900 4956
rect 4676 4946 4900 4951
rect 4666 4890 4676 4946
rect 4732 4900 4900 4946
rect 4956 4900 4966 4956
rect 5450 4900 5460 4956
rect 5516 4900 5684 4956
rect 5740 4900 5750 4956
rect 6346 4900 6356 4956
rect 6412 4900 7812 4956
rect 7868 4951 7951 4956
rect 8250 4951 8372 4956
rect 7868 4900 8372 4951
rect 8428 4900 8438 4956
rect 12954 4900 12964 4956
rect 13020 4905 13412 4956
rect 13468 4905 13478 4961
rect 13020 4900 13468 4905
rect 13626 4900 13636 4956
rect 13692 4900 14980 4956
rect 15036 4900 15764 4956
rect 15820 4900 15830 4956
rect 18106 4900 18116 4956
rect 18172 4900 18340 4956
rect 18396 4900 18406 4956
rect 19226 4900 19236 4956
rect 19292 4900 21476 4956
rect 21532 4900 23044 4956
rect 23100 4900 23110 4956
rect 23706 4900 23716 4956
rect 23772 4900 24108 4956
rect 4732 4895 4843 4900
rect 7883 4895 8307 4900
rect 4732 4890 4742 4895
rect 2090 4788 2100 4844
rect 2156 4788 2884 4844
rect 2940 4834 4127 4844
rect 2940 4788 5012 4834
rect 4062 4778 5012 4788
rect 5068 4778 5078 4834
rect 6234 4788 6244 4844
rect 6300 4788 7252 4844
rect 7308 4788 7318 4844
rect 11946 4788 11956 4844
rect 12012 4824 22932 4844
rect 12012 4788 13412 4824
rect 13402 4768 13412 4788
rect 13468 4788 22932 4824
rect 22988 4788 22998 4844
rect 13468 4768 13478 4788
rect 1754 4676 1764 4732
rect 1820 4676 2212 4732
rect 2268 4722 4012 4732
rect 2268 4676 5124 4722
rect 3949 4666 5124 4676
rect 5180 4666 5190 4722
rect 5898 4676 5908 4732
rect 5964 4676 8484 4732
rect 8540 4676 8550 4732
rect 1866 4564 1876 4620
rect 1932 4564 3780 4620
rect 3836 4564 3846 4620
rect 16408 4508 16460 4564
rect 16516 4508 16616 4564
rect 16672 4508 16772 4564
rect 16828 4508 16928 4564
rect 16984 4508 17084 4564
rect 17140 4508 17192 4564
rect 1306 4452 1316 4508
rect 1372 4452 4004 4508
rect 4060 4452 4900 4508
rect 4956 4452 4966 4508
rect 298 4340 308 4396
rect 364 4340 756 4396
rect 812 4340 2884 4396
rect 2940 4340 4228 4396
rect 4284 4340 4294 4396
rect 9930 4340 9940 4396
rect 9996 4340 10836 4396
rect 10892 4340 12404 4396
rect 12460 4340 13300 4396
rect 13356 4340 13366 4396
rect 1530 4228 1540 4284
rect 1596 4228 2772 4284
rect 2828 4228 3668 4284
rect 3724 4264 4900 4284
rect 3724 4228 4116 4264
rect 4106 4208 4116 4228
rect 4172 4228 4900 4264
rect 4956 4228 6916 4284
rect 6972 4228 6982 4284
rect 13850 4228 13860 4284
rect 13916 4228 16996 4284
rect 17052 4228 17062 4284
rect 4172 4208 4182 4228
rect 410 4116 420 4172
rect 476 4116 980 4172
rect 1036 4116 1046 4172
rect 1642 4116 1652 4172
rect 1708 4116 2324 4172
rect 2380 4116 3892 4172
rect 3948 4116 3958 4172
rect 4554 4116 4564 4172
rect 4620 4116 5236 4172
rect 5292 4116 5684 4172
rect 5740 4116 5750 4172
rect 7354 4116 7364 4172
rect 7420 4116 8820 4172
rect 8876 4116 8886 4172
rect 12730 4116 12740 4172
rect 12796 4116 14308 4172
rect 14364 4116 14374 4172
rect 14970 4116 14980 4172
rect 15036 4116 17444 4172
rect 17500 4116 19012 4172
rect 19068 4116 19078 4172
rect 10169 4060 10225 4070
rect 2202 4004 2212 4060
rect 2268 4004 2660 4060
rect 2716 4004 2726 4060
rect 3098 4004 3108 4060
rect 3164 4004 4452 4060
rect 4508 4004 4564 4060
rect 4620 4004 4630 4060
rect 7578 4004 7588 4060
rect 7644 4004 10047 4060
rect 10103 4004 10113 4060
rect 10225 4004 10500 4060
rect 10556 4004 10566 4060
rect 15082 4004 15092 4060
rect 15148 4040 17296 4060
rect 15148 4035 17500 4040
rect 15148 4004 17444 4035
rect 10169 3994 10225 4004
rect 17221 3984 17444 4004
rect 17434 3979 17444 3984
rect 17500 3979 17510 4035
rect 18890 4004 18900 4060
rect 18956 4004 19908 4060
rect 19964 4004 19974 4060
rect 22810 4004 22820 4060
rect 22876 4004 24108 4060
rect 1978 3892 1988 3948
rect 2044 3892 3780 3948
rect 3836 3892 3846 3948
rect 8474 3780 8484 3836
rect 8540 3780 8820 3836
rect 8876 3780 8886 3836
rect 15530 3780 15540 3836
rect 15596 3780 17220 3836
rect 17276 3780 18228 3836
rect 18284 3780 20020 3836
rect 20076 3780 20086 3836
rect 5992 3612 6044 3668
rect 6100 3612 6200 3668
rect 6256 3612 6356 3668
rect 6412 3612 6512 3668
rect 6568 3612 6668 3668
rect 6724 3612 6776 3668
rect 17770 3556 17780 3612
rect 17836 3556 20244 3612
rect 20300 3556 20310 3612
rect 5236 3444 8260 3500
rect 8316 3444 8326 3500
rect 5236 3388 5292 3444
rect 8708 3398 8764 3500
rect 16202 3444 16212 3500
rect 16268 3444 18340 3500
rect 18396 3444 18406 3500
rect 2538 3332 2548 3388
rect 2604 3332 4116 3388
rect 4172 3332 5236 3388
rect 5292 3332 5302 3388
rect 5786 3332 5796 3388
rect 5852 3332 8036 3388
rect 8092 3332 8102 3388
rect 8698 3342 8708 3398
rect 8764 3342 8774 3398
rect 10042 3337 10052 3393
rect 10108 3388 10118 3393
rect 10108 3337 10276 3388
rect 10052 3332 10276 3337
rect 10332 3332 10342 3388
rect 15978 3332 15988 3388
rect 16044 3332 17220 3388
rect 17276 3332 17286 3388
rect 19002 3332 19012 3388
rect 19068 3332 20804 3388
rect 20860 3332 20870 3388
rect 21802 3337 21812 3393
rect 21868 3388 21878 3393
rect 21868 3337 22596 3388
rect 21812 3332 22596 3337
rect 22652 3332 22662 3388
rect 23034 3332 23044 3388
rect 23100 3332 24108 3388
rect 858 3220 868 3276
rect 924 3220 1316 3276
rect 1372 3220 1382 3276
rect 1530 3220 1540 3276
rect 1596 3220 1876 3276
rect 1932 3220 1942 3276
rect 2202 3220 2212 3276
rect 2268 3220 3444 3276
rect 3500 3220 3510 3276
rect 7354 3220 7364 3276
rect 7420 3220 8932 3276
rect 8988 3220 8998 3276
rect 10052 3271 12516 3276
rect 10042 3215 10052 3271
rect 10108 3220 12516 3271
rect 12572 3220 12582 3276
rect 14746 3240 14756 3296
rect 14812 3276 14822 3296
rect 14812 3240 16996 3276
rect 14756 3220 16996 3240
rect 17052 3220 17062 3276
rect 19338 3220 19348 3276
rect 19404 3220 21588 3276
rect 21644 3220 21654 3276
rect 21914 3220 21924 3276
rect 21980 3220 23380 3276
rect 23436 3220 23446 3276
rect 10108 3215 10118 3220
rect 23380 3164 23436 3220
rect 2538 3108 2548 3164
rect 2604 3108 2996 3164
rect 3052 3108 3780 3164
rect 3836 3108 5012 3164
rect 5068 3108 5078 3164
rect 7354 3108 7364 3164
rect 7420 3108 7476 3164
rect 7532 3108 7542 3164
rect 7914 3108 7924 3164
rect 7980 3108 8708 3164
rect 8764 3108 8774 3164
rect 11498 3108 11508 3164
rect 11564 3108 12832 3164
rect 12888 3108 12898 3164
rect 12959 3108 12969 3164
rect 13025 3108 13188 3164
rect 13244 3108 13254 3164
rect 14186 3108 14196 3164
rect 14252 3108 14644 3164
rect 14700 3108 15316 3164
rect 15372 3108 15382 3164
rect 16090 3108 16100 3164
rect 16156 3108 17892 3164
rect 17948 3108 17958 3164
rect 18666 3108 18676 3164
rect 18732 3108 22596 3164
rect 22652 3108 22662 3164
rect 23380 3108 24108 3164
rect 298 2996 308 3052
rect 364 2996 644 3052
rect 700 2996 710 3052
rect 4218 2996 4228 3052
rect 4284 2996 5460 3052
rect 5516 3032 7259 3052
rect 5516 3027 7532 3032
rect 5516 2996 7476 3027
rect 7203 2976 7476 2996
rect 7466 2971 7476 2976
rect 7532 2971 7542 3027
rect 10378 2996 10388 3052
rect 10444 2996 14084 3052
rect 14140 2996 14756 3052
rect 14812 2996 14822 3052
rect 3882 2884 3892 2940
rect 3948 2884 4788 2940
rect 4844 2884 4854 2940
rect 12282 2884 12292 2940
rect 12348 2884 12964 2940
rect 13020 2884 13030 2940
rect 3546 2772 3556 2828
rect 3612 2772 4228 2828
rect 4284 2772 4294 2828
rect 1866 2716 1876 2721
rect 1642 2660 1652 2716
rect 1708 2665 1876 2716
rect 1932 2665 1942 2721
rect 4440 2719 4452 2775
rect 4508 2719 4676 2775
rect 4732 2719 4742 2775
rect 16408 2716 16460 2772
rect 16516 2716 16616 2772
rect 16672 2716 16772 2772
rect 16828 2716 16928 2772
rect 16984 2716 17084 2772
rect 17140 2716 17192 2772
rect 1708 2660 1932 2665
rect 18442 2660 18452 2716
rect 18508 2660 22484 2716
rect 22540 2660 22550 2716
rect 1876 2599 2100 2604
rect 1866 2543 1876 2599
rect 1932 2548 2100 2599
rect 2156 2548 2166 2604
rect 1932 2543 1942 2548
rect 7364 2492 7420 2604
rect 12170 2548 12180 2604
rect 12236 2548 16212 2604
rect 16268 2548 16772 2604
rect 16828 2548 16838 2604
rect 17098 2548 17108 2604
rect 17164 2548 17780 2604
rect 17836 2548 17846 2604
rect 17994 2548 18004 2604
rect 18060 2548 18788 2604
rect 18844 2548 18854 2604
rect 7354 2436 7364 2492
rect 7420 2436 7430 2492
rect 7690 2441 7700 2497
rect 7756 2492 7766 2497
rect 7756 2441 8708 2492
rect 7700 2436 8708 2441
rect 8764 2436 8774 2492
rect 13290 2436 13300 2492
rect 13356 2436 14420 2492
rect 14476 2436 16324 2492
rect 16380 2436 16390 2492
rect 18330 2436 18340 2492
rect 18396 2436 20580 2492
rect 20636 2436 20646 2492
rect 5562 2324 5572 2380
rect 5628 2375 7756 2380
rect 5628 2324 7700 2375
rect 7690 2319 7700 2324
rect 7756 2319 7766 2375
rect 8586 2324 8596 2380
rect 8652 2324 8820 2380
rect 8876 2324 9940 2380
rect 9996 2324 11732 2380
rect 11788 2324 11798 2380
rect 12282 2324 12292 2380
rect 12348 2324 14532 2380
rect 14588 2324 14598 2380
rect 14848 2324 14858 2380
rect 14914 2324 15316 2380
rect 15372 2324 15856 2380
rect 15912 2324 15922 2380
rect 15983 2324 15993 2380
rect 16049 2324 16548 2380
rect 16604 2324 17556 2380
rect 17612 2324 17622 2380
rect 18554 2324 18564 2380
rect 18620 2324 18788 2380
rect 18844 2324 18854 2380
rect 5002 2212 5012 2268
rect 5068 2212 6244 2268
rect 6300 2258 7457 2268
rect 6300 2253 8036 2258
rect 6300 2212 7588 2253
rect 7397 2202 7588 2212
rect 7578 2197 7588 2202
rect 7644 2202 8036 2253
rect 8092 2202 8102 2258
rect 8250 2217 8260 2273
rect 8316 2268 8326 2273
rect 8316 2217 9268 2268
rect 8260 2212 9268 2217
rect 9324 2212 9334 2268
rect 10490 2212 10500 2268
rect 10556 2212 11060 2268
rect 11116 2212 11126 2268
rect 12058 2212 12068 2268
rect 12124 2212 14420 2268
rect 14476 2212 14644 2268
rect 14700 2212 14710 2268
rect 14766 2212 14776 2268
rect 14832 2212 18452 2268
rect 18508 2212 18518 2268
rect 7644 2197 7654 2202
rect 4218 2100 4228 2156
rect 4284 2100 4676 2156
rect 4732 2100 5348 2156
rect 5404 2100 5414 2156
rect 9594 2100 9604 2156
rect 9660 2100 10164 2156
rect 10220 2100 10612 2156
rect 10668 2100 10678 2156
rect 14522 2100 14532 2156
rect 14588 2100 17668 2156
rect 17724 2100 17734 2156
rect 10378 1988 10388 2044
rect 10444 1988 11172 2044
rect 11228 1988 11238 2044
rect 13626 1988 13636 2044
rect 13692 1988 15647 2044
rect 15703 1988 15713 2044
rect 15774 1988 15784 2044
rect 15840 1988 18116 2044
rect 18172 1988 18182 2044
rect 5992 1820 6044 1876
rect 6100 1820 6200 1876
rect 6256 1820 6356 1876
rect 6412 1820 6512 1876
rect 6568 1820 6668 1876
rect 6724 1820 6776 1876
rect 1754 1652 1764 1708
rect 1820 1652 3668 1708
rect 3724 1652 3734 1708
rect 13962 1652 13972 1708
rect 14028 1652 15204 1708
rect 15260 1652 15270 1708
rect 16762 1652 16772 1708
rect 16828 1652 17556 1708
rect 17612 1652 17622 1708
rect 10490 1596 10500 1601
rect 1418 1540 1428 1596
rect 1484 1540 2324 1596
rect 2380 1540 3556 1596
rect 3612 1540 7700 1596
rect 7756 1540 8484 1596
rect 8540 1540 9940 1596
rect 9996 1545 10500 1596
rect 10556 1545 10566 1601
rect 9996 1540 10556 1545
rect 13514 1540 13524 1596
rect 13580 1540 14756 1596
rect 14812 1540 14822 1596
rect 18218 1540 18228 1596
rect 18284 1540 22260 1596
rect 22316 1540 22326 1596
rect 13402 1484 13412 1489
rect 2426 1428 2436 1484
rect 2492 1428 4004 1484
rect 4060 1428 4070 1484
rect 4890 1428 4900 1484
rect 4956 1428 6020 1484
rect 6076 1428 8596 1484
rect 8652 1428 8662 1484
rect 10490 1408 10500 1484
rect 10556 1433 13412 1484
rect 13468 1433 13478 1489
rect 10556 1428 13468 1433
rect 15306 1428 15316 1484
rect 15372 1479 16156 1484
rect 15372 1428 16212 1479
rect 10556 1408 10566 1428
rect 16091 1423 16212 1428
rect 16268 1423 16436 1479
rect 16492 1423 16502 1479
rect 17882 1428 17892 1484
rect 17948 1428 18004 1484
rect 18060 1428 18070 1484
rect 18554 1428 18564 1484
rect 18620 1428 20244 1484
rect 20300 1428 20310 1484
rect 20458 1428 20468 1484
rect 20524 1428 22372 1484
rect 22428 1428 22438 1484
rect 1194 1316 1204 1372
rect 1260 1316 2772 1372
rect 2828 1316 2838 1372
rect 3658 1316 3668 1372
rect 3724 1316 4340 1372
rect 4396 1316 4406 1372
rect 6346 1316 6356 1372
rect 6412 1316 7140 1372
rect 7196 1316 8148 1372
rect 8204 1316 9828 1372
rect 9884 1316 9894 1372
rect 12618 1316 12628 1372
rect 12684 1316 14532 1372
rect 14588 1316 14598 1372
rect 16584 1367 18228 1372
rect 15978 1311 15988 1367
rect 16044 1316 18228 1367
rect 18284 1316 18294 1372
rect 21130 1316 21140 1372
rect 21196 1316 21588 1372
rect 21644 1316 21654 1372
rect 23706 1316 23716 1372
rect 23772 1316 24108 1372
rect 16044 1311 16641 1316
rect 8698 1204 8708 1260
rect 8764 1204 12292 1260
rect 12348 1204 12358 1260
rect 15194 1204 15204 1260
rect 15260 1204 15540 1260
rect 15596 1204 15606 1260
rect 17546 1204 17556 1260
rect 17612 1204 18340 1260
rect 18396 1204 20356 1260
rect 20412 1204 20422 1260
rect 1642 980 1652 1036
rect 1708 980 8260 1036
rect 8316 980 8326 1036
rect 8708 924 8764 1036
rect 16408 924 16460 980
rect 16516 924 16616 980
rect 16672 924 16772 980
rect 16828 924 16928 980
rect 16984 924 17084 980
rect 17140 924 17192 980
rect 3098 868 3108 924
rect 3164 868 8708 924
rect 8764 868 8774 924
rect 15082 868 15092 924
rect 15148 868 15540 924
rect 15596 868 15606 924
rect 858 756 868 812
rect 924 756 11508 812
rect 11564 756 12740 812
rect 12796 756 14980 812
rect 15036 756 15876 812
rect 15932 756 15942 812
rect 17658 756 17668 812
rect 17724 756 18788 812
rect 18844 756 18854 812
rect 4666 644 4676 700
rect 4732 644 5684 700
rect 5740 644 9268 700
rect 9324 644 10388 700
rect 10444 644 10454 700
rect 12282 644 12292 700
rect 12348 644 13412 700
rect 13468 644 14084 700
rect 14140 644 14150 700
rect 15082 644 15092 700
rect 15148 644 15540 700
rect 15596 644 15606 700
rect 17322 644 17332 700
rect 17388 644 18900 700
rect 18956 644 18966 700
rect 3882 532 3892 588
rect 3948 532 4900 588
rect 4956 532 4966 588
rect 7588 476 7644 588
rect 11386 532 11396 588
rect 11452 532 12852 588
rect 12908 532 13524 588
rect 13580 532 13748 588
rect 13804 532 13814 588
rect 14522 532 14532 588
rect 14588 532 15204 588
rect 15260 532 15270 588
rect 16650 532 16660 588
rect 16716 532 17556 588
rect 17612 532 17622 588
rect 18330 532 18340 588
rect 18396 532 20692 588
rect 20748 532 20758 588
rect 1866 420 1876 476
rect 1932 420 7588 476
rect 7644 420 7654 476
rect 22484 420 22596 476
rect 22652 420 22662 476
rect 18330 84 18340 140
rect 18396 84 19124 140
rect 19180 84 19190 140
rect 5992 28 6044 84
rect 6100 28 6200 84
rect 6256 28 6356 84
rect 6412 28 6512 84
rect 6568 28 6668 84
rect 6724 28 6776 84
<< via3 >>
rect 16460 20636 16516 20692
rect 16616 20636 16672 20692
rect 16772 20636 16828 20692
rect 16928 20636 16984 20692
rect 17084 20636 17140 20692
rect 6044 19740 6100 19796
rect 6200 19740 6256 19796
rect 6356 19740 6412 19796
rect 6512 19740 6568 19796
rect 6668 19740 6724 19796
rect 23716 19684 23772 19740
rect 4788 19256 4844 19292
rect 4788 19236 4844 19256
rect 4788 18900 4844 18956
rect 16460 18844 16516 18900
rect 16616 18844 16672 18900
rect 16772 18844 16828 18900
rect 16928 18844 16984 18900
rect 17084 18844 17140 18900
rect 22372 18452 22428 18508
rect 308 18228 364 18284
rect 10948 18228 11004 18284
rect 3108 18024 3164 18060
rect 3108 18004 3164 18024
rect 6044 17948 6100 18004
rect 6200 17948 6256 18004
rect 6356 17948 6412 18004
rect 6512 17948 6568 18004
rect 6668 17948 6724 18004
rect 23716 17332 23772 17388
rect 10164 17220 10220 17276
rect 16460 17052 16516 17108
rect 16616 17052 16672 17108
rect 16772 17052 16828 17108
rect 16928 17052 16984 17108
rect 17084 17052 17140 17108
rect 2548 16996 2604 17052
rect 308 16884 364 16940
rect 2548 16533 2604 16589
rect 10948 16436 11004 16492
rect 6044 16156 6100 16212
rect 6200 16156 6256 16212
rect 6356 16156 6412 16212
rect 6512 16156 6568 16212
rect 6668 16156 6724 16212
rect 23716 15764 23772 15820
rect 16460 15260 16516 15316
rect 16616 15260 16672 15316
rect 16772 15260 16828 15316
rect 16928 15260 16984 15316
rect 17084 15260 17140 15316
rect 21028 15092 21084 15148
rect 6044 14364 6100 14420
rect 6200 14364 6256 14420
rect 6356 14364 6412 14420
rect 6512 14364 6568 14420
rect 6668 14364 6724 14420
rect 14420 14084 14476 14140
rect 3108 13860 3164 13916
rect 13636 13524 13692 13580
rect 16460 13468 16516 13524
rect 16616 13468 16672 13524
rect 16772 13468 16828 13524
rect 16928 13468 16984 13524
rect 17084 13468 17140 13524
rect 11732 13076 11788 13132
rect 17668 12852 17724 12908
rect 1428 12740 1484 12796
rect 6044 12572 6100 12628
rect 6200 12572 6256 12628
rect 6356 12572 6412 12628
rect 6512 12572 6568 12628
rect 6668 12572 6724 12628
rect 20020 11956 20076 12012
rect 22372 11956 22428 12012
rect 16460 11676 16516 11732
rect 16616 11676 16672 11732
rect 16772 11676 16828 11732
rect 16928 11676 16984 11732
rect 17084 11676 17140 11732
rect 1428 11396 1484 11452
rect 14980 10948 15036 11004
rect 6044 10780 6100 10836
rect 6200 10780 6256 10836
rect 6356 10780 6412 10836
rect 6512 10780 6568 10836
rect 6668 10780 6724 10836
rect 2548 10388 2604 10444
rect 18564 10388 18620 10444
rect 11732 10164 11788 10220
rect 16460 9884 16516 9940
rect 16616 9884 16672 9940
rect 16772 9884 16828 9940
rect 16928 9884 16984 9940
rect 17084 9884 17140 9940
rect 15204 9738 15260 9794
rect 15428 9626 15484 9682
rect 21252 9604 21308 9660
rect 6044 8988 6100 9044
rect 6200 8988 6256 9044
rect 6356 8988 6412 9044
rect 6512 8988 6568 9044
rect 6668 8988 6724 9044
rect 17912 8820 17968 8876
rect 17668 8708 17724 8764
rect 4340 8596 4396 8652
rect 11620 8596 11676 8652
rect 23716 8596 23772 8652
rect 9044 8484 9100 8540
rect 14420 8484 14476 8540
rect 5460 8260 5516 8316
rect 16460 8092 16516 8148
rect 16616 8092 16672 8148
rect 16772 8092 16828 8148
rect 16928 8092 16984 8148
rect 17084 8092 17140 8148
rect 15204 7924 15260 7980
rect 17332 7924 17388 7980
rect 21028 7812 21084 7868
rect 17332 7700 17388 7756
rect 4900 7476 4956 7532
rect 6044 7196 6100 7252
rect 6200 7196 6256 7252
rect 6356 7196 6412 7252
rect 6512 7196 6568 7252
rect 6668 7196 6724 7252
rect 14980 6804 15036 6860
rect 15428 6804 15484 6860
rect 20020 6692 20076 6748
rect 17332 6468 17388 6524
rect 16460 6300 16516 6356
rect 16616 6300 16672 6356
rect 16772 6300 16828 6356
rect 16928 6300 16984 6356
rect 17084 6300 17140 6356
rect 9044 6020 9100 6076
rect 18004 5796 18060 5852
rect 18788 5796 18844 5852
rect 21252 5796 21308 5852
rect 3780 5572 3836 5628
rect 4335 5460 4391 5516
rect 6044 5404 6100 5460
rect 6200 5404 6256 5460
rect 6356 5404 6412 5460
rect 6512 5404 6568 5460
rect 6668 5404 6724 5460
rect 5460 5348 5516 5404
rect 13636 5348 13692 5404
rect 4564 5012 4620 5068
rect 15535 5022 15591 5073
rect 15535 5017 15591 5022
rect 4900 4900 4956 4956
rect 18340 4900 18396 4956
rect 16460 4508 16516 4564
rect 16616 4508 16672 4564
rect 16772 4508 16828 4564
rect 16928 4508 16984 4564
rect 17084 4508 17140 4564
rect 4564 4004 4620 4060
rect 7588 4004 7644 4060
rect 10169 4004 10225 4060
rect 10500 4004 10556 4060
rect 6044 3612 6100 3668
rect 6200 3612 6256 3668
rect 6356 3612 6412 3668
rect 6512 3612 6568 3668
rect 6668 3612 6724 3668
rect 8708 3342 8764 3398
rect 22596 3332 22652 3388
rect 3780 3108 3836 3164
rect 7364 3108 7420 3164
rect 16460 2716 16516 2772
rect 16616 2716 16672 2772
rect 16772 2716 16828 2772
rect 16928 2716 16984 2772
rect 17084 2716 17140 2772
rect 7364 2436 7420 2492
rect 18564 2324 18620 2380
rect 6044 1820 6100 1876
rect 6200 1820 6256 1876
rect 6356 1820 6412 1876
rect 6512 1820 6568 1876
rect 6668 1820 6724 1876
rect 10500 1464 10556 1484
rect 10500 1428 10556 1464
rect 18004 1428 18060 1484
rect 18340 1204 18396 1260
rect 16460 924 16516 980
rect 16616 924 16672 980
rect 16772 924 16828 980
rect 16928 924 16984 980
rect 17084 924 17140 980
rect 8708 868 8764 924
rect 18788 756 18844 812
rect 15540 644 15596 700
rect 7588 420 7644 476
rect 22596 420 22652 476
rect 6044 28 6100 84
rect 6200 28 6256 84
rect 6356 28 6412 84
rect 6512 28 6568 84
rect 6668 28 6724 84
<< metal4 >>
rect 16408 20702 17192 20718
rect 16408 20626 16441 20702
rect 16517 20692 16655 20702
rect 16731 20692 16869 20702
rect 16945 20692 17083 20702
rect 16517 20636 16616 20692
rect 16731 20636 16772 20692
rect 16828 20636 16869 20692
rect 16984 20636 17083 20692
rect 16517 20626 16655 20636
rect 16731 20626 16869 20636
rect 16945 20626 17083 20636
rect 17159 20626 17192 20702
rect 16408 20610 17192 20626
rect 5992 19806 6776 19822
rect 5992 19730 6025 19806
rect 6101 19796 6239 19806
rect 6315 19796 6453 19806
rect 6529 19796 6667 19806
rect 6101 19740 6200 19796
rect 6315 19740 6356 19796
rect 6412 19740 6453 19796
rect 6568 19740 6667 19796
rect 6101 19730 6239 19740
rect 6315 19730 6453 19740
rect 6529 19730 6667 19740
rect 6743 19730 6776 19806
rect 5992 19714 6776 19730
rect 23716 19740 23772 19750
rect 4788 19292 4844 19302
rect 4788 18956 4844 19236
rect 4788 18890 4844 18900
rect 16408 18910 17192 18926
rect 16408 18834 16441 18910
rect 16517 18900 16655 18910
rect 16731 18900 16869 18910
rect 16945 18900 17083 18910
rect 16517 18844 16616 18900
rect 16731 18844 16772 18900
rect 16828 18844 16869 18900
rect 16984 18844 17083 18900
rect 16517 18834 16655 18844
rect 16731 18834 16869 18844
rect 16945 18834 17083 18844
rect 17159 18834 17192 18910
rect 16408 18818 17192 18834
rect 22372 18508 22428 18518
rect 308 18284 364 18294
rect 308 16940 364 18228
rect 10948 18284 11004 18294
rect 3108 18060 3164 18070
rect 308 16874 364 16884
rect 2548 17052 2604 17062
rect 2548 16589 2604 16996
rect 1428 12796 1484 12806
rect 1428 11452 1484 12740
rect 1428 11386 1484 11396
rect 2548 10444 2604 16533
rect 3108 13916 3164 18004
rect 5992 18014 6776 18030
rect 5992 17938 6025 18014
rect 6101 18004 6239 18014
rect 6315 18004 6453 18014
rect 6529 18004 6667 18014
rect 6101 17948 6200 18004
rect 6315 17948 6356 18004
rect 6412 17948 6453 18004
rect 6568 17948 6667 18004
rect 6101 17938 6239 17948
rect 6315 17938 6453 17948
rect 6529 17938 6667 17948
rect 6743 17938 6776 18014
rect 5992 17922 6776 17938
rect 10164 17276 10220 17286
rect 5992 16222 6776 16238
rect 5992 16146 6025 16222
rect 6101 16212 6239 16222
rect 6315 16212 6453 16222
rect 6529 16212 6667 16222
rect 6101 16156 6200 16212
rect 6315 16156 6356 16212
rect 6412 16156 6453 16212
rect 6568 16156 6667 16212
rect 6101 16146 6239 16156
rect 6315 16146 6453 16156
rect 6529 16146 6667 16156
rect 6743 16146 6776 16222
rect 5992 16130 6776 16146
rect 5992 14430 6776 14446
rect 5992 14354 6025 14430
rect 6101 14420 6239 14430
rect 6315 14420 6453 14430
rect 6529 14420 6667 14430
rect 6101 14364 6200 14420
rect 6315 14364 6356 14420
rect 6412 14364 6453 14420
rect 6568 14364 6667 14420
rect 6101 14354 6239 14364
rect 6315 14354 6453 14364
rect 6529 14354 6667 14364
rect 6743 14354 6776 14430
rect 5992 14338 6776 14354
rect 3108 13850 3164 13860
rect 5992 12638 6776 12654
rect 5992 12562 6025 12638
rect 6101 12628 6239 12638
rect 6315 12628 6453 12638
rect 6529 12628 6667 12638
rect 6101 12572 6200 12628
rect 6315 12572 6356 12628
rect 6412 12572 6453 12628
rect 6568 12572 6667 12628
rect 6101 12562 6239 12572
rect 6315 12562 6453 12572
rect 6529 12562 6667 12572
rect 6743 12562 6776 12638
rect 5992 12546 6776 12562
rect 5992 10846 6776 10862
rect 5992 10770 6025 10846
rect 6101 10836 6239 10846
rect 6315 10836 6453 10846
rect 6529 10836 6667 10846
rect 6101 10780 6200 10836
rect 6315 10780 6356 10836
rect 6412 10780 6453 10836
rect 6568 10780 6667 10836
rect 6101 10770 6239 10780
rect 6315 10770 6453 10780
rect 6529 10770 6667 10780
rect 6743 10770 6776 10846
rect 5992 10754 6776 10770
rect 2548 10378 2604 10388
rect 5992 9054 6776 9070
rect 5992 8978 6025 9054
rect 6101 9044 6239 9054
rect 6315 9044 6453 9054
rect 6529 9044 6667 9054
rect 6101 8988 6200 9044
rect 6315 8988 6356 9044
rect 6412 8988 6453 9044
rect 6568 8988 6667 9044
rect 6101 8978 6239 8988
rect 6315 8978 6453 8988
rect 6529 8978 6667 8988
rect 6743 8978 6776 9054
rect 5992 8962 6776 8978
rect 4340 8652 4396 8662
rect 3780 5628 3836 5638
rect 3780 3164 3836 5572
rect 4340 5526 4396 8596
rect 9044 8540 9100 8550
rect 5460 8316 5516 8326
rect 4335 5516 4396 5526
rect 4391 5460 4396 5516
rect 4900 7532 4956 7542
rect 4335 5450 4391 5460
rect 4564 5068 4620 5078
rect 4564 4060 4620 5012
rect 4900 4956 4956 7476
rect 5460 5404 5516 8260
rect 5992 7262 6776 7278
rect 5992 7186 6025 7262
rect 6101 7252 6239 7262
rect 6315 7252 6453 7262
rect 6529 7252 6667 7262
rect 6101 7196 6200 7252
rect 6315 7196 6356 7252
rect 6412 7196 6453 7252
rect 6568 7196 6667 7252
rect 6101 7186 6239 7196
rect 6315 7186 6453 7196
rect 6529 7186 6667 7196
rect 6743 7186 6776 7262
rect 5992 7170 6776 7186
rect 9044 6076 9100 8484
rect 9044 6010 9100 6020
rect 5992 5470 6776 5486
rect 5992 5394 6025 5470
rect 6101 5460 6239 5470
rect 6315 5460 6453 5470
rect 6529 5460 6667 5470
rect 6101 5404 6200 5460
rect 6315 5404 6356 5460
rect 6412 5404 6453 5460
rect 6568 5404 6667 5460
rect 6101 5394 6239 5404
rect 6315 5394 6453 5404
rect 6529 5394 6667 5404
rect 6743 5394 6776 5470
rect 5992 5378 6776 5394
rect 5460 5338 5516 5348
rect 4900 4890 4956 4900
rect 10164 4070 10220 17220
rect 10948 16492 11004 18228
rect 16408 17118 17192 17134
rect 16408 17042 16441 17118
rect 16517 17108 16655 17118
rect 16731 17108 16869 17118
rect 16945 17108 17083 17118
rect 16517 17052 16616 17108
rect 16731 17052 16772 17108
rect 16828 17052 16869 17108
rect 16984 17052 17083 17108
rect 16517 17042 16655 17052
rect 16731 17042 16869 17052
rect 16945 17042 17083 17052
rect 17159 17042 17192 17118
rect 16408 17026 17192 17042
rect 10948 16426 11004 16436
rect 16408 15326 17192 15342
rect 16408 15250 16441 15326
rect 16517 15316 16655 15326
rect 16731 15316 16869 15326
rect 16945 15316 17083 15326
rect 16517 15260 16616 15316
rect 16731 15260 16772 15316
rect 16828 15260 16869 15316
rect 16984 15260 17083 15316
rect 16517 15250 16655 15260
rect 16731 15250 16869 15260
rect 16945 15250 17083 15260
rect 17159 15250 17192 15326
rect 16408 15234 17192 15250
rect 21028 15148 21084 15158
rect 14420 14140 14476 14150
rect 13636 13580 13692 13590
rect 11732 13132 11788 13142
rect 11732 10220 11788 13076
rect 11732 10154 11788 10164
rect 11610 8886 11686 8896
rect 11610 8800 11686 8810
rect 11620 8652 11676 8800
rect 11620 8586 11676 8596
rect 13636 5404 13692 13524
rect 14420 8540 14476 14084
rect 16408 13534 17192 13550
rect 16408 13458 16441 13534
rect 16517 13524 16655 13534
rect 16731 13524 16869 13534
rect 16945 13524 17083 13534
rect 16517 13468 16616 13524
rect 16731 13468 16772 13524
rect 16828 13468 16869 13524
rect 16984 13468 17083 13524
rect 16517 13458 16655 13468
rect 16731 13458 16869 13468
rect 16945 13458 17083 13468
rect 17159 13458 17192 13534
rect 16408 13442 17192 13458
rect 17668 12908 17724 12918
rect 16408 11742 17192 11758
rect 16408 11666 16441 11742
rect 16517 11732 16655 11742
rect 16731 11732 16869 11742
rect 16945 11732 17083 11742
rect 16517 11676 16616 11732
rect 16731 11676 16772 11732
rect 16828 11676 16869 11732
rect 16984 11676 17083 11732
rect 16517 11666 16655 11676
rect 16731 11666 16869 11676
rect 16945 11666 17083 11676
rect 17159 11666 17192 11742
rect 16408 11650 17192 11666
rect 14420 8474 14476 8484
rect 14980 11004 15036 11014
rect 14980 6860 15036 10948
rect 16408 9950 17192 9966
rect 16408 9874 16441 9950
rect 16517 9940 16655 9950
rect 16731 9940 16869 9950
rect 16945 9940 17083 9950
rect 16517 9884 16616 9940
rect 16731 9884 16772 9940
rect 16828 9884 16869 9940
rect 16984 9884 17083 9940
rect 16517 9874 16655 9884
rect 16731 9874 16869 9884
rect 16945 9874 17083 9884
rect 17159 9874 17192 9950
rect 16408 9858 17192 9874
rect 15204 9794 15260 9804
rect 15204 7980 15260 9738
rect 15204 7914 15260 7924
rect 15428 9682 15484 9692
rect 14980 6794 15036 6804
rect 15428 6860 15484 9626
rect 17668 8764 17724 12852
rect 20020 12012 20076 12022
rect 18564 10444 18620 10454
rect 17882 8886 17958 8896
rect 17958 8876 17968 8886
rect 17968 8820 18060 8876
rect 17958 8810 17968 8820
rect 17882 8800 17958 8810
rect 17668 8698 17724 8708
rect 16408 8158 17192 8174
rect 16408 8082 16441 8158
rect 16517 8148 16655 8158
rect 16731 8148 16869 8158
rect 16945 8148 17083 8158
rect 16517 8092 16616 8148
rect 16731 8092 16772 8148
rect 16828 8092 16869 8148
rect 16984 8092 17083 8148
rect 16517 8082 16655 8092
rect 16731 8082 16869 8092
rect 16945 8082 17083 8092
rect 17159 8082 17192 8158
rect 16408 8066 17192 8082
rect 15428 6794 15484 6804
rect 17332 7980 17388 7990
rect 17332 7756 17388 7924
rect 17332 6524 17388 7700
rect 17332 6458 17388 6468
rect 16408 6366 17192 6382
rect 16408 6290 16441 6366
rect 16517 6356 16655 6366
rect 16731 6356 16869 6366
rect 16945 6356 17083 6366
rect 16517 6300 16616 6356
rect 16731 6300 16772 6356
rect 16828 6300 16869 6356
rect 16984 6300 17083 6356
rect 16517 6290 16655 6300
rect 16731 6290 16869 6300
rect 16945 6290 17083 6300
rect 17159 6290 17192 6366
rect 16408 6274 17192 6290
rect 13636 5338 13692 5348
rect 18004 5852 18060 5862
rect 15535 5073 15591 5083
rect 15591 5017 15596 5073
rect 15535 5007 15596 5017
rect 4564 3994 4620 4004
rect 7588 4060 7644 4070
rect 10164 4060 10225 4070
rect 10164 4004 10169 4060
rect 5992 3678 6776 3694
rect 5992 3602 6025 3678
rect 6101 3668 6239 3678
rect 6315 3668 6453 3678
rect 6529 3668 6667 3678
rect 6101 3612 6200 3668
rect 6315 3612 6356 3668
rect 6412 3612 6453 3668
rect 6568 3612 6667 3668
rect 6101 3602 6239 3612
rect 6315 3602 6453 3612
rect 6529 3602 6667 3612
rect 6743 3602 6776 3678
rect 5992 3586 6776 3602
rect 3780 3098 3836 3108
rect 7364 3164 7420 3174
rect 7364 2492 7420 3108
rect 7364 2426 7420 2436
rect 5992 1886 6776 1902
rect 5992 1810 6025 1886
rect 6101 1876 6239 1886
rect 6315 1876 6453 1886
rect 6529 1876 6667 1886
rect 6101 1820 6200 1876
rect 6315 1820 6356 1876
rect 6412 1820 6453 1876
rect 6568 1820 6667 1876
rect 6101 1810 6239 1820
rect 6315 1810 6453 1820
rect 6529 1810 6667 1820
rect 6743 1810 6776 1886
rect 5992 1794 6776 1810
rect 7588 476 7644 4004
rect 10169 3994 10225 4004
rect 10500 4060 10556 4070
rect 8708 3398 8764 3408
rect 8708 924 8764 3342
rect 10500 1484 10556 4004
rect 10500 1418 10556 1428
rect 8708 858 8764 868
rect 15540 700 15596 5007
rect 16408 4574 17192 4590
rect 16408 4498 16441 4574
rect 16517 4564 16655 4574
rect 16731 4564 16869 4574
rect 16945 4564 17083 4574
rect 16517 4508 16616 4564
rect 16731 4508 16772 4564
rect 16828 4508 16869 4564
rect 16984 4508 17083 4564
rect 16517 4498 16655 4508
rect 16731 4498 16869 4508
rect 16945 4498 17083 4508
rect 17159 4498 17192 4574
rect 16408 4482 17192 4498
rect 16408 2782 17192 2798
rect 16408 2706 16441 2782
rect 16517 2772 16655 2782
rect 16731 2772 16869 2782
rect 16945 2772 17083 2782
rect 16517 2716 16616 2772
rect 16731 2716 16772 2772
rect 16828 2716 16869 2772
rect 16984 2716 17083 2772
rect 16517 2706 16655 2716
rect 16731 2706 16869 2716
rect 16945 2706 17083 2716
rect 17159 2706 17192 2782
rect 16408 2690 17192 2706
rect 18004 1484 18060 5796
rect 18004 1418 18060 1428
rect 18340 4956 18396 4966
rect 18340 1260 18396 4900
rect 18564 2380 18620 10388
rect 20020 6748 20076 11956
rect 21028 7868 21084 15092
rect 22372 12012 22428 18452
rect 23716 17388 23772 19684
rect 23716 17322 23772 17332
rect 22372 11946 22428 11956
rect 23716 15820 23772 15830
rect 21028 7802 21084 7812
rect 21252 9660 21308 9670
rect 20020 6682 20076 6692
rect 18564 2314 18620 2324
rect 18788 5852 18844 5862
rect 18340 1194 18396 1204
rect 16408 990 17192 1006
rect 16408 914 16441 990
rect 16517 980 16655 990
rect 16731 980 16869 990
rect 16945 980 17083 990
rect 16517 924 16616 980
rect 16731 924 16772 980
rect 16828 924 16869 980
rect 16984 924 17083 980
rect 16517 914 16655 924
rect 16731 914 16869 924
rect 16945 914 17083 924
rect 17159 914 17192 990
rect 16408 898 17192 914
rect 18788 812 18844 5796
rect 21252 5852 21308 9604
rect 23716 8652 23772 15764
rect 23716 8586 23772 8596
rect 21252 5786 21308 5796
rect 18788 746 18844 756
rect 22596 3388 22652 3398
rect 15540 634 15596 644
rect 7588 410 7644 420
rect 22596 476 22652 3332
rect 22596 410 22652 420
rect 5992 94 6776 110
rect 5992 18 6025 94
rect 6101 84 6239 94
rect 6315 84 6453 94
rect 6529 84 6667 94
rect 6101 28 6200 84
rect 6315 28 6356 84
rect 6412 28 6453 84
rect 6568 28 6667 84
rect 6101 18 6239 28
rect 6315 18 6453 28
rect 6529 18 6667 28
rect 6743 18 6776 94
rect 5992 2 6776 18
<< viatp >>
rect 16441 20692 16517 20702
rect 16655 20692 16731 20702
rect 16869 20692 16945 20702
rect 17083 20692 17159 20702
rect 16441 20636 16460 20692
rect 16460 20636 16516 20692
rect 16516 20636 16517 20692
rect 16655 20636 16672 20692
rect 16672 20636 16731 20692
rect 16869 20636 16928 20692
rect 16928 20636 16945 20692
rect 17083 20636 17084 20692
rect 17084 20636 17140 20692
rect 17140 20636 17159 20692
rect 16441 20626 16517 20636
rect 16655 20626 16731 20636
rect 16869 20626 16945 20636
rect 17083 20626 17159 20636
rect 6025 19796 6101 19806
rect 6239 19796 6315 19806
rect 6453 19796 6529 19806
rect 6667 19796 6743 19806
rect 6025 19740 6044 19796
rect 6044 19740 6100 19796
rect 6100 19740 6101 19796
rect 6239 19740 6256 19796
rect 6256 19740 6315 19796
rect 6453 19740 6512 19796
rect 6512 19740 6529 19796
rect 6667 19740 6668 19796
rect 6668 19740 6724 19796
rect 6724 19740 6743 19796
rect 6025 19730 6101 19740
rect 6239 19730 6315 19740
rect 6453 19730 6529 19740
rect 6667 19730 6743 19740
rect 16441 18900 16517 18910
rect 16655 18900 16731 18910
rect 16869 18900 16945 18910
rect 17083 18900 17159 18910
rect 16441 18844 16460 18900
rect 16460 18844 16516 18900
rect 16516 18844 16517 18900
rect 16655 18844 16672 18900
rect 16672 18844 16731 18900
rect 16869 18844 16928 18900
rect 16928 18844 16945 18900
rect 17083 18844 17084 18900
rect 17084 18844 17140 18900
rect 17140 18844 17159 18900
rect 16441 18834 16517 18844
rect 16655 18834 16731 18844
rect 16869 18834 16945 18844
rect 17083 18834 17159 18844
rect 6025 18004 6101 18014
rect 6239 18004 6315 18014
rect 6453 18004 6529 18014
rect 6667 18004 6743 18014
rect 6025 17948 6044 18004
rect 6044 17948 6100 18004
rect 6100 17948 6101 18004
rect 6239 17948 6256 18004
rect 6256 17948 6315 18004
rect 6453 17948 6512 18004
rect 6512 17948 6529 18004
rect 6667 17948 6668 18004
rect 6668 17948 6724 18004
rect 6724 17948 6743 18004
rect 6025 17938 6101 17948
rect 6239 17938 6315 17948
rect 6453 17938 6529 17948
rect 6667 17938 6743 17948
rect 6025 16212 6101 16222
rect 6239 16212 6315 16222
rect 6453 16212 6529 16222
rect 6667 16212 6743 16222
rect 6025 16156 6044 16212
rect 6044 16156 6100 16212
rect 6100 16156 6101 16212
rect 6239 16156 6256 16212
rect 6256 16156 6315 16212
rect 6453 16156 6512 16212
rect 6512 16156 6529 16212
rect 6667 16156 6668 16212
rect 6668 16156 6724 16212
rect 6724 16156 6743 16212
rect 6025 16146 6101 16156
rect 6239 16146 6315 16156
rect 6453 16146 6529 16156
rect 6667 16146 6743 16156
rect 6025 14420 6101 14430
rect 6239 14420 6315 14430
rect 6453 14420 6529 14430
rect 6667 14420 6743 14430
rect 6025 14364 6044 14420
rect 6044 14364 6100 14420
rect 6100 14364 6101 14420
rect 6239 14364 6256 14420
rect 6256 14364 6315 14420
rect 6453 14364 6512 14420
rect 6512 14364 6529 14420
rect 6667 14364 6668 14420
rect 6668 14364 6724 14420
rect 6724 14364 6743 14420
rect 6025 14354 6101 14364
rect 6239 14354 6315 14364
rect 6453 14354 6529 14364
rect 6667 14354 6743 14364
rect 6025 12628 6101 12638
rect 6239 12628 6315 12638
rect 6453 12628 6529 12638
rect 6667 12628 6743 12638
rect 6025 12572 6044 12628
rect 6044 12572 6100 12628
rect 6100 12572 6101 12628
rect 6239 12572 6256 12628
rect 6256 12572 6315 12628
rect 6453 12572 6512 12628
rect 6512 12572 6529 12628
rect 6667 12572 6668 12628
rect 6668 12572 6724 12628
rect 6724 12572 6743 12628
rect 6025 12562 6101 12572
rect 6239 12562 6315 12572
rect 6453 12562 6529 12572
rect 6667 12562 6743 12572
rect 6025 10836 6101 10846
rect 6239 10836 6315 10846
rect 6453 10836 6529 10846
rect 6667 10836 6743 10846
rect 6025 10780 6044 10836
rect 6044 10780 6100 10836
rect 6100 10780 6101 10836
rect 6239 10780 6256 10836
rect 6256 10780 6315 10836
rect 6453 10780 6512 10836
rect 6512 10780 6529 10836
rect 6667 10780 6668 10836
rect 6668 10780 6724 10836
rect 6724 10780 6743 10836
rect 6025 10770 6101 10780
rect 6239 10770 6315 10780
rect 6453 10770 6529 10780
rect 6667 10770 6743 10780
rect 6025 9044 6101 9054
rect 6239 9044 6315 9054
rect 6453 9044 6529 9054
rect 6667 9044 6743 9054
rect 6025 8988 6044 9044
rect 6044 8988 6100 9044
rect 6100 8988 6101 9044
rect 6239 8988 6256 9044
rect 6256 8988 6315 9044
rect 6453 8988 6512 9044
rect 6512 8988 6529 9044
rect 6667 8988 6668 9044
rect 6668 8988 6724 9044
rect 6724 8988 6743 9044
rect 6025 8978 6101 8988
rect 6239 8978 6315 8988
rect 6453 8978 6529 8988
rect 6667 8978 6743 8988
rect 6025 7252 6101 7262
rect 6239 7252 6315 7262
rect 6453 7252 6529 7262
rect 6667 7252 6743 7262
rect 6025 7196 6044 7252
rect 6044 7196 6100 7252
rect 6100 7196 6101 7252
rect 6239 7196 6256 7252
rect 6256 7196 6315 7252
rect 6453 7196 6512 7252
rect 6512 7196 6529 7252
rect 6667 7196 6668 7252
rect 6668 7196 6724 7252
rect 6724 7196 6743 7252
rect 6025 7186 6101 7196
rect 6239 7186 6315 7196
rect 6453 7186 6529 7196
rect 6667 7186 6743 7196
rect 6025 5460 6101 5470
rect 6239 5460 6315 5470
rect 6453 5460 6529 5470
rect 6667 5460 6743 5470
rect 6025 5404 6044 5460
rect 6044 5404 6100 5460
rect 6100 5404 6101 5460
rect 6239 5404 6256 5460
rect 6256 5404 6315 5460
rect 6453 5404 6512 5460
rect 6512 5404 6529 5460
rect 6667 5404 6668 5460
rect 6668 5404 6724 5460
rect 6724 5404 6743 5460
rect 6025 5394 6101 5404
rect 6239 5394 6315 5404
rect 6453 5394 6529 5404
rect 6667 5394 6743 5404
rect 16441 17108 16517 17118
rect 16655 17108 16731 17118
rect 16869 17108 16945 17118
rect 17083 17108 17159 17118
rect 16441 17052 16460 17108
rect 16460 17052 16516 17108
rect 16516 17052 16517 17108
rect 16655 17052 16672 17108
rect 16672 17052 16731 17108
rect 16869 17052 16928 17108
rect 16928 17052 16945 17108
rect 17083 17052 17084 17108
rect 17084 17052 17140 17108
rect 17140 17052 17159 17108
rect 16441 17042 16517 17052
rect 16655 17042 16731 17052
rect 16869 17042 16945 17052
rect 17083 17042 17159 17052
rect 16441 15316 16517 15326
rect 16655 15316 16731 15326
rect 16869 15316 16945 15326
rect 17083 15316 17159 15326
rect 16441 15260 16460 15316
rect 16460 15260 16516 15316
rect 16516 15260 16517 15316
rect 16655 15260 16672 15316
rect 16672 15260 16731 15316
rect 16869 15260 16928 15316
rect 16928 15260 16945 15316
rect 17083 15260 17084 15316
rect 17084 15260 17140 15316
rect 17140 15260 17159 15316
rect 16441 15250 16517 15260
rect 16655 15250 16731 15260
rect 16869 15250 16945 15260
rect 17083 15250 17159 15260
rect 11610 8810 11686 8886
rect 16441 13524 16517 13534
rect 16655 13524 16731 13534
rect 16869 13524 16945 13534
rect 17083 13524 17159 13534
rect 16441 13468 16460 13524
rect 16460 13468 16516 13524
rect 16516 13468 16517 13524
rect 16655 13468 16672 13524
rect 16672 13468 16731 13524
rect 16869 13468 16928 13524
rect 16928 13468 16945 13524
rect 17083 13468 17084 13524
rect 17084 13468 17140 13524
rect 17140 13468 17159 13524
rect 16441 13458 16517 13468
rect 16655 13458 16731 13468
rect 16869 13458 16945 13468
rect 17083 13458 17159 13468
rect 16441 11732 16517 11742
rect 16655 11732 16731 11742
rect 16869 11732 16945 11742
rect 17083 11732 17159 11742
rect 16441 11676 16460 11732
rect 16460 11676 16516 11732
rect 16516 11676 16517 11732
rect 16655 11676 16672 11732
rect 16672 11676 16731 11732
rect 16869 11676 16928 11732
rect 16928 11676 16945 11732
rect 17083 11676 17084 11732
rect 17084 11676 17140 11732
rect 17140 11676 17159 11732
rect 16441 11666 16517 11676
rect 16655 11666 16731 11676
rect 16869 11666 16945 11676
rect 17083 11666 17159 11676
rect 16441 9940 16517 9950
rect 16655 9940 16731 9950
rect 16869 9940 16945 9950
rect 17083 9940 17159 9950
rect 16441 9884 16460 9940
rect 16460 9884 16516 9940
rect 16516 9884 16517 9940
rect 16655 9884 16672 9940
rect 16672 9884 16731 9940
rect 16869 9884 16928 9940
rect 16928 9884 16945 9940
rect 17083 9884 17084 9940
rect 17084 9884 17140 9940
rect 17140 9884 17159 9940
rect 16441 9874 16517 9884
rect 16655 9874 16731 9884
rect 16869 9874 16945 9884
rect 17083 9874 17159 9884
rect 17882 8876 17958 8886
rect 17882 8820 17912 8876
rect 17912 8820 17958 8876
rect 17882 8810 17958 8820
rect 16441 8148 16517 8158
rect 16655 8148 16731 8158
rect 16869 8148 16945 8158
rect 17083 8148 17159 8158
rect 16441 8092 16460 8148
rect 16460 8092 16516 8148
rect 16516 8092 16517 8148
rect 16655 8092 16672 8148
rect 16672 8092 16731 8148
rect 16869 8092 16928 8148
rect 16928 8092 16945 8148
rect 17083 8092 17084 8148
rect 17084 8092 17140 8148
rect 17140 8092 17159 8148
rect 16441 8082 16517 8092
rect 16655 8082 16731 8092
rect 16869 8082 16945 8092
rect 17083 8082 17159 8092
rect 16441 6356 16517 6366
rect 16655 6356 16731 6366
rect 16869 6356 16945 6366
rect 17083 6356 17159 6366
rect 16441 6300 16460 6356
rect 16460 6300 16516 6356
rect 16516 6300 16517 6356
rect 16655 6300 16672 6356
rect 16672 6300 16731 6356
rect 16869 6300 16928 6356
rect 16928 6300 16945 6356
rect 17083 6300 17084 6356
rect 17084 6300 17140 6356
rect 17140 6300 17159 6356
rect 16441 6290 16517 6300
rect 16655 6290 16731 6300
rect 16869 6290 16945 6300
rect 17083 6290 17159 6300
rect 6025 3668 6101 3678
rect 6239 3668 6315 3678
rect 6453 3668 6529 3678
rect 6667 3668 6743 3678
rect 6025 3612 6044 3668
rect 6044 3612 6100 3668
rect 6100 3612 6101 3668
rect 6239 3612 6256 3668
rect 6256 3612 6315 3668
rect 6453 3612 6512 3668
rect 6512 3612 6529 3668
rect 6667 3612 6668 3668
rect 6668 3612 6724 3668
rect 6724 3612 6743 3668
rect 6025 3602 6101 3612
rect 6239 3602 6315 3612
rect 6453 3602 6529 3612
rect 6667 3602 6743 3612
rect 6025 1876 6101 1886
rect 6239 1876 6315 1886
rect 6453 1876 6529 1886
rect 6667 1876 6743 1886
rect 6025 1820 6044 1876
rect 6044 1820 6100 1876
rect 6100 1820 6101 1876
rect 6239 1820 6256 1876
rect 6256 1820 6315 1876
rect 6453 1820 6512 1876
rect 6512 1820 6529 1876
rect 6667 1820 6668 1876
rect 6668 1820 6724 1876
rect 6724 1820 6743 1876
rect 6025 1810 6101 1820
rect 6239 1810 6315 1820
rect 6453 1810 6529 1820
rect 6667 1810 6743 1820
rect 16441 4564 16517 4574
rect 16655 4564 16731 4574
rect 16869 4564 16945 4574
rect 17083 4564 17159 4574
rect 16441 4508 16460 4564
rect 16460 4508 16516 4564
rect 16516 4508 16517 4564
rect 16655 4508 16672 4564
rect 16672 4508 16731 4564
rect 16869 4508 16928 4564
rect 16928 4508 16945 4564
rect 17083 4508 17084 4564
rect 17084 4508 17140 4564
rect 17140 4508 17159 4564
rect 16441 4498 16517 4508
rect 16655 4498 16731 4508
rect 16869 4498 16945 4508
rect 17083 4498 17159 4508
rect 16441 2772 16517 2782
rect 16655 2772 16731 2782
rect 16869 2772 16945 2782
rect 17083 2772 17159 2782
rect 16441 2716 16460 2772
rect 16460 2716 16516 2772
rect 16516 2716 16517 2772
rect 16655 2716 16672 2772
rect 16672 2716 16731 2772
rect 16869 2716 16928 2772
rect 16928 2716 16945 2772
rect 17083 2716 17084 2772
rect 17084 2716 17140 2772
rect 17140 2716 17159 2772
rect 16441 2706 16517 2716
rect 16655 2706 16731 2716
rect 16869 2706 16945 2716
rect 17083 2706 17159 2716
rect 16441 980 16517 990
rect 16655 980 16731 990
rect 16869 980 16945 990
rect 17083 980 17159 990
rect 16441 924 16460 980
rect 16460 924 16516 980
rect 16516 924 16517 980
rect 16655 924 16672 980
rect 16672 924 16731 980
rect 16869 924 16928 980
rect 16928 924 16945 980
rect 17083 924 17084 980
rect 17084 924 17140 980
rect 17140 924 17159 980
rect 16441 914 16517 924
rect 16655 914 16731 924
rect 16869 914 16945 924
rect 17083 914 17159 924
rect 6025 84 6101 94
rect 6239 84 6315 94
rect 6453 84 6529 94
rect 6667 84 6743 94
rect 6025 28 6044 84
rect 6044 28 6100 84
rect 6100 28 6101 84
rect 6239 28 6256 84
rect 6256 28 6315 84
rect 6453 28 6512 84
rect 6512 28 6529 84
rect 6667 28 6668 84
rect 6668 28 6724 84
rect 6724 28 6743 84
rect 6025 18 6101 28
rect 6239 18 6315 28
rect 6453 18 6529 28
rect 6667 18 6743 28
<< metaltp >>
rect 16408 20702 16500 20814
rect 17100 20702 17192 20814
rect 16408 20626 16441 20702
rect 17159 20626 17192 20702
rect 16408 20514 16500 20626
rect 17100 20514 17192 20626
rect 5992 19806 6084 19918
rect 6684 19806 6776 19918
rect 5992 19730 6025 19806
rect 6743 19730 6776 19806
rect 5992 19618 6084 19730
rect 6684 19618 6776 19730
rect 16408 18910 16500 19022
rect 17100 18910 17192 19022
rect 16408 18834 16441 18910
rect 17159 18834 17192 18910
rect 16408 18722 16500 18834
rect 17100 18722 17192 18834
rect 5992 18014 6084 18126
rect 6684 18014 6776 18126
rect 5992 17938 6025 18014
rect 6743 17938 6776 18014
rect 5992 17826 6084 17938
rect 6684 17826 6776 17938
rect 16408 17118 16500 17230
rect 17100 17118 17192 17230
rect 16408 17042 16441 17118
rect 17159 17042 17192 17118
rect 16408 16930 16500 17042
rect 17100 16930 17192 17042
rect 5992 16222 6084 16334
rect 6684 16222 6776 16334
rect 5992 16146 6025 16222
rect 6743 16146 6776 16222
rect 5992 16034 6084 16146
rect 6684 16034 6776 16146
rect 16408 15326 16500 15438
rect 17100 15326 17192 15438
rect 16408 15250 16441 15326
rect 17159 15250 17192 15326
rect 16408 15138 16500 15250
rect 17100 15138 17192 15250
rect 5992 14430 6084 14542
rect 6684 14430 6776 14542
rect 5992 14354 6025 14430
rect 6743 14354 6776 14430
rect 5992 14242 6084 14354
rect 6684 14242 6776 14354
rect 16408 13534 16500 13646
rect 17100 13534 17192 13646
rect 16408 13458 16441 13534
rect 17159 13458 17192 13534
rect 16408 13346 16500 13458
rect 17100 13346 17192 13458
rect 5992 12638 6084 12750
rect 6684 12638 6776 12750
rect 5992 12562 6025 12638
rect 6743 12562 6776 12638
rect 5992 12450 6084 12562
rect 6684 12450 6776 12562
rect 16408 11742 16500 11854
rect 17100 11742 17192 11854
rect 16408 11666 16441 11742
rect 17159 11666 17192 11742
rect 16408 11554 16500 11666
rect 17100 11554 17192 11666
rect 5992 10846 6084 10958
rect 6684 10846 6776 10958
rect 5992 10770 6025 10846
rect 6743 10770 6776 10846
rect 5992 10658 6084 10770
rect 6684 10658 6776 10770
rect 16408 9950 16500 10062
rect 17100 9950 17192 10062
rect 16408 9874 16441 9950
rect 17159 9874 17192 9950
rect 16408 9762 16500 9874
rect 17100 9762 17192 9874
rect 5992 9054 6084 9166
rect 6684 9054 6776 9166
rect 5992 8978 6025 9054
rect 6743 8978 6776 9054
rect 5992 8866 6084 8978
rect 6684 8866 6776 8978
rect 11594 8892 11702 8902
rect 17866 8892 17974 8902
rect 11594 8886 17974 8892
rect 11594 8810 11610 8886
rect 11686 8810 17882 8886
rect 17958 8810 17974 8886
rect 11594 8804 17974 8810
rect 11594 8794 11702 8804
rect 17866 8794 17974 8804
rect 16408 8158 16500 8270
rect 17100 8158 17192 8270
rect 16408 8082 16441 8158
rect 17159 8082 17192 8158
rect 16408 7970 16500 8082
rect 17100 7970 17192 8082
rect 5992 7262 6084 7374
rect 6684 7262 6776 7374
rect 5992 7186 6025 7262
rect 6743 7186 6776 7262
rect 5992 7074 6084 7186
rect 6684 7074 6776 7186
rect 16408 6366 16500 6478
rect 17100 6366 17192 6478
rect 16408 6290 16441 6366
rect 17159 6290 17192 6366
rect 16408 6178 16500 6290
rect 17100 6178 17192 6290
rect 5992 5470 6084 5582
rect 6684 5470 6776 5582
rect 5992 5394 6025 5470
rect 6743 5394 6776 5470
rect 5992 5282 6084 5394
rect 6684 5282 6776 5394
rect 16408 4574 16500 4686
rect 17100 4574 17192 4686
rect 16408 4498 16441 4574
rect 17159 4498 17192 4574
rect 16408 4386 16500 4498
rect 17100 4386 17192 4498
rect 5992 3678 6084 3790
rect 6684 3678 6776 3790
rect 5992 3602 6025 3678
rect 6743 3602 6776 3678
rect 5992 3490 6084 3602
rect 6684 3490 6776 3602
rect 16408 2782 16500 2894
rect 17100 2782 17192 2894
rect 16408 2706 16441 2782
rect 17159 2706 17192 2782
rect 16408 2594 16500 2706
rect 17100 2594 17192 2706
rect 5992 1886 6084 1998
rect 6684 1886 6776 1998
rect 5992 1810 6025 1886
rect 6743 1810 6776 1886
rect 5992 1698 6084 1810
rect 6684 1698 6776 1810
rect 16408 990 16500 1102
rect 17100 990 17192 1102
rect 16408 914 16441 990
rect 17159 914 17192 990
rect 16408 802 16500 914
rect 17100 802 17192 914
rect 5992 94 6084 206
rect 6684 94 6776 206
rect 5992 18 6025 94
rect 6743 18 6776 94
rect 5992 -94 6084 18
rect 6684 -94 6776 18
<< viatpl >>
rect 16500 20702 17100 20814
rect 16500 20626 16517 20702
rect 16517 20626 16655 20702
rect 16655 20626 16731 20702
rect 16731 20626 16869 20702
rect 16869 20626 16945 20702
rect 16945 20626 17083 20702
rect 17083 20626 17100 20702
rect 16500 20514 17100 20626
rect 6084 19806 6684 19918
rect 6084 19730 6101 19806
rect 6101 19730 6239 19806
rect 6239 19730 6315 19806
rect 6315 19730 6453 19806
rect 6453 19730 6529 19806
rect 6529 19730 6667 19806
rect 6667 19730 6684 19806
rect 6084 19618 6684 19730
rect 16500 18910 17100 19022
rect 16500 18834 16517 18910
rect 16517 18834 16655 18910
rect 16655 18834 16731 18910
rect 16731 18834 16869 18910
rect 16869 18834 16945 18910
rect 16945 18834 17083 18910
rect 17083 18834 17100 18910
rect 16500 18722 17100 18834
rect 6084 18014 6684 18126
rect 6084 17938 6101 18014
rect 6101 17938 6239 18014
rect 6239 17938 6315 18014
rect 6315 17938 6453 18014
rect 6453 17938 6529 18014
rect 6529 17938 6667 18014
rect 6667 17938 6684 18014
rect 6084 17826 6684 17938
rect 16500 17118 17100 17230
rect 16500 17042 16517 17118
rect 16517 17042 16655 17118
rect 16655 17042 16731 17118
rect 16731 17042 16869 17118
rect 16869 17042 16945 17118
rect 16945 17042 17083 17118
rect 17083 17042 17100 17118
rect 16500 16930 17100 17042
rect 6084 16222 6684 16334
rect 6084 16146 6101 16222
rect 6101 16146 6239 16222
rect 6239 16146 6315 16222
rect 6315 16146 6453 16222
rect 6453 16146 6529 16222
rect 6529 16146 6667 16222
rect 6667 16146 6684 16222
rect 6084 16034 6684 16146
rect 16500 15326 17100 15438
rect 16500 15250 16517 15326
rect 16517 15250 16655 15326
rect 16655 15250 16731 15326
rect 16731 15250 16869 15326
rect 16869 15250 16945 15326
rect 16945 15250 17083 15326
rect 17083 15250 17100 15326
rect 16500 15138 17100 15250
rect 6084 14430 6684 14542
rect 6084 14354 6101 14430
rect 6101 14354 6239 14430
rect 6239 14354 6315 14430
rect 6315 14354 6453 14430
rect 6453 14354 6529 14430
rect 6529 14354 6667 14430
rect 6667 14354 6684 14430
rect 6084 14242 6684 14354
rect 16500 13534 17100 13646
rect 16500 13458 16517 13534
rect 16517 13458 16655 13534
rect 16655 13458 16731 13534
rect 16731 13458 16869 13534
rect 16869 13458 16945 13534
rect 16945 13458 17083 13534
rect 17083 13458 17100 13534
rect 16500 13346 17100 13458
rect 6084 12638 6684 12750
rect 6084 12562 6101 12638
rect 6101 12562 6239 12638
rect 6239 12562 6315 12638
rect 6315 12562 6453 12638
rect 6453 12562 6529 12638
rect 6529 12562 6667 12638
rect 6667 12562 6684 12638
rect 6084 12450 6684 12562
rect 16500 11742 17100 11854
rect 16500 11666 16517 11742
rect 16517 11666 16655 11742
rect 16655 11666 16731 11742
rect 16731 11666 16869 11742
rect 16869 11666 16945 11742
rect 16945 11666 17083 11742
rect 17083 11666 17100 11742
rect 16500 11554 17100 11666
rect 6084 10846 6684 10958
rect 6084 10770 6101 10846
rect 6101 10770 6239 10846
rect 6239 10770 6315 10846
rect 6315 10770 6453 10846
rect 6453 10770 6529 10846
rect 6529 10770 6667 10846
rect 6667 10770 6684 10846
rect 6084 10658 6684 10770
rect 16500 9950 17100 10062
rect 16500 9874 16517 9950
rect 16517 9874 16655 9950
rect 16655 9874 16731 9950
rect 16731 9874 16869 9950
rect 16869 9874 16945 9950
rect 16945 9874 17083 9950
rect 17083 9874 17100 9950
rect 16500 9762 17100 9874
rect 6084 9054 6684 9166
rect 6084 8978 6101 9054
rect 6101 8978 6239 9054
rect 6239 8978 6315 9054
rect 6315 8978 6453 9054
rect 6453 8978 6529 9054
rect 6529 8978 6667 9054
rect 6667 8978 6684 9054
rect 6084 8866 6684 8978
rect 16500 8158 17100 8270
rect 16500 8082 16517 8158
rect 16517 8082 16655 8158
rect 16655 8082 16731 8158
rect 16731 8082 16869 8158
rect 16869 8082 16945 8158
rect 16945 8082 17083 8158
rect 17083 8082 17100 8158
rect 16500 7970 17100 8082
rect 6084 7262 6684 7374
rect 6084 7186 6101 7262
rect 6101 7186 6239 7262
rect 6239 7186 6315 7262
rect 6315 7186 6453 7262
rect 6453 7186 6529 7262
rect 6529 7186 6667 7262
rect 6667 7186 6684 7262
rect 6084 7074 6684 7186
rect 16500 6366 17100 6478
rect 16500 6290 16517 6366
rect 16517 6290 16655 6366
rect 16655 6290 16731 6366
rect 16731 6290 16869 6366
rect 16869 6290 16945 6366
rect 16945 6290 17083 6366
rect 17083 6290 17100 6366
rect 16500 6178 17100 6290
rect 6084 5470 6684 5582
rect 6084 5394 6101 5470
rect 6101 5394 6239 5470
rect 6239 5394 6315 5470
rect 6315 5394 6453 5470
rect 6453 5394 6529 5470
rect 6529 5394 6667 5470
rect 6667 5394 6684 5470
rect 6084 5282 6684 5394
rect 16500 4574 17100 4686
rect 16500 4498 16517 4574
rect 16517 4498 16655 4574
rect 16655 4498 16731 4574
rect 16731 4498 16869 4574
rect 16869 4498 16945 4574
rect 16945 4498 17083 4574
rect 17083 4498 17100 4574
rect 16500 4386 17100 4498
rect 6084 3678 6684 3790
rect 6084 3602 6101 3678
rect 6101 3602 6239 3678
rect 6239 3602 6315 3678
rect 6315 3602 6453 3678
rect 6453 3602 6529 3678
rect 6529 3602 6667 3678
rect 6667 3602 6684 3678
rect 6084 3490 6684 3602
rect 16500 2782 17100 2894
rect 16500 2706 16517 2782
rect 16517 2706 16655 2782
rect 16655 2706 16731 2782
rect 16731 2706 16869 2782
rect 16869 2706 16945 2782
rect 16945 2706 17083 2782
rect 17083 2706 17100 2782
rect 16500 2594 17100 2706
rect 6084 1886 6684 1998
rect 6084 1810 6101 1886
rect 6101 1810 6239 1886
rect 6239 1810 6315 1886
rect 6315 1810 6453 1886
rect 6453 1810 6529 1886
rect 6529 1810 6667 1886
rect 6667 1810 6684 1886
rect 6084 1698 6684 1810
rect 16500 990 17100 1102
rect 16500 914 16517 990
rect 16517 914 16655 990
rect 16655 914 16731 990
rect 16731 914 16869 990
rect 16869 914 16945 990
rect 16945 914 17083 990
rect 17083 914 17100 990
rect 16500 802 17100 914
rect 6084 94 6684 206
rect 6084 18 6101 94
rect 6101 18 6239 94
rect 6239 18 6315 94
rect 6315 18 6453 94
rect 6453 18 6529 94
rect 6529 18 6667 94
rect 6667 18 6684 94
rect 6084 -94 6684 18
<< metaltpl >>
rect 5992 19918 6776 20944
rect 5992 19618 6084 19918
rect 6684 19618 6776 19918
rect 5992 18126 6776 19618
rect 5992 17826 6084 18126
rect 6684 17826 6776 18126
rect 5992 16334 6776 17826
rect 5992 16034 6084 16334
rect 6684 16034 6776 16334
rect 5992 14542 6776 16034
rect 5992 14242 6084 14542
rect 6684 14242 6776 14542
rect 5992 12750 6776 14242
rect 5992 12450 6084 12750
rect 6684 12450 6776 12750
rect 5992 10958 6776 12450
rect 5992 10658 6084 10958
rect 6684 10658 6776 10958
rect 5992 9166 6776 10658
rect 5992 8866 6084 9166
rect 6684 8866 6776 9166
rect 5992 7374 6776 8866
rect 5992 7074 6084 7374
rect 6684 7074 6776 7374
rect 5992 5582 6776 7074
rect 5992 5282 6084 5582
rect 6684 5282 6776 5582
rect 5992 3790 6776 5282
rect 5992 3490 6084 3790
rect 6684 3490 6776 3790
rect 5992 1998 6776 3490
rect 5992 1698 6084 1998
rect 6684 1698 6776 1998
rect 5992 206 6776 1698
rect 5992 -94 6084 206
rect 6684 -94 6776 206
rect 5992 -336 6776 -94
rect 16408 20814 17192 20944
rect 16408 20514 16500 20814
rect 17100 20514 17192 20814
rect 16408 19022 17192 20514
rect 16408 18722 16500 19022
rect 17100 18722 17192 19022
rect 16408 17230 17192 18722
rect 16408 16930 16500 17230
rect 17100 16930 17192 17230
rect 16408 15438 17192 16930
rect 16408 15138 16500 15438
rect 17100 15138 17192 15438
rect 16408 13646 17192 15138
rect 16408 13346 16500 13646
rect 17100 13346 17192 13646
rect 16408 11854 17192 13346
rect 16408 11554 16500 11854
rect 17100 11554 17192 11854
rect 16408 10062 17192 11554
rect 16408 9762 16500 10062
rect 17100 9762 17192 10062
rect 16408 8270 17192 9762
rect 16408 7970 16500 8270
rect 17100 7970 17192 8270
rect 16408 6478 17192 7970
rect 16408 6178 16500 6478
rect 17100 6178 17192 6478
rect 16408 4686 17192 6178
rect 16408 4386 16500 4686
rect 17100 4386 17192 4686
rect 16408 2894 17192 4386
rect 16408 2594 16500 2894
rect 17100 2594 17192 2894
rect 16408 1102 17192 2594
rect 16408 802 16500 1102
rect 17100 802 17192 1102
rect 16408 -336 17192 802
use DFRRQ_3VX4  DFRRQ_3VX4_32 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 56 0 -1 20664
box 0 0 3584 896
use NA2_3VX0  NA2_3VX0_19 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 4088 0 -1 20664
box 0 0 448 896
use NA3_3VX0  NA3_3VX0_19 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 4648 0 -1 20664
box 0 0 560 896
use NA3I2_3VX1  NA3I2_3VX1_4 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 4648 0 -1 20664
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_NA2_3VX0_16 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 5432 0 -1 20664
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_16
timestamp 1529525674
transform 1 0 5992 0 -1 20664
box 0 0 448 896
use DECAP7_3V  DECAP7_3V_22_0_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 6440 0 -1 20664
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_33
timestamp 1529525674
transform 1 0 7224 0 -1 20664
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_33
timestamp 1529525674
transform 1 0 7784 0 -1 20664
box 0 0 3584 896
use DECAP5_3V  DECAP5_3V_0_MU2_3VX0_4
timestamp 1529525674
transform -1 0 11928 0 -1 20664
box 0 0 560 896
use MU2_3VX0  MU2_3VX0_4 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 13048 0 -1 20664
box 0 0 1120 896
use MU2_3VX0  MU2_3VX0_7
timestamp 1529525674
transform 1 0 13272 0 -1 20664
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_36
timestamp 1529525674
transform 1 0 14392 0 -1 20664
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_22_1_0
timestamp 1529525674
transform 1 0 14952 0 -1 20664
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_36
timestamp 1529525674
transform 1 0 15736 0 -1 20664
box 0 0 3584 896
use BU_3VX2  BU_3VX2_31 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 19320 0 -1 20664
box 0 0 672 896
use LOGIC0_3V  LOGIC0_3V_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 19992 0 -1 20664
box 0 0 560 896
use DECAP5_3V  DECAP5_3V_0_BU_3VX2_17
timestamp 1529525674
transform 1 0 20552 0 -1 20664
box 0 0 560 896
use BU_3VX2  BU_3VX2_17
timestamp 1529525674
transform 1 0 21112 0 -1 20664
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_DFRSQ_3VX4_6
timestamp 1529525674
transform 1 0 280 0 1 18872
box 0 0 560 896
use DFRSQ_3VX4  DFRSQ_3VX4_6 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 840 0 1 18872
box 0 0 3360 896
use NA3_3VX0  NA3_3VX0_20
timestamp 1529525674
transform -1 0 4760 0 1 18872
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_17
timestamp 1529525674
transform -1 0 5208 0 1 18872
box 0 0 448 896
use IN_3VX0  IN_3VX0_21 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 5544 0 1 18872
box 0 0 336 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_31
timestamp 1529525674
transform -1 0 6104 0 1 18872
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_21_0_0
timestamp 1529525674
transform -1 0 6888 0 1 18872
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_31
timestamp 1529525674
transform -1 0 10472 0 1 18872
box 0 0 3584 896
use DECAP5_3V  DECAP5_3V_0_DFFSQ_3VX1_1
timestamp 1529525674
transform -1 0 11032 0 1 18872
box 0 0 560 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_7 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 13048 0 -1 20664
box 0 -80 224 976
use DFFSQ_3VX1  DFFSQ_3VX1_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 13832 0 1 18872
box 0 0 2800 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_15
timestamp 1529525674
transform 1 0 13832 0 1 18872
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_15
timestamp 1529525674
transform 1 0 14392 0 1 18872
box 0 0 3584 896
use DECAP7_3V  DECAP7_3V_21_1_0
timestamp 1529525674
transform 1 0 17976 0 1 18872
box 0 0 784 896
use AND2_3VX0  AND2_3VX0_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 18760 0 1 18872
box 0 0 672 896
use AND2_3VX0  AND2_3VX0_3
timestamp 1529525674
transform 1 0 19432 0 1 18872
box 0 0 672 896
use BU_3VX2  BU_3VX2_32
timestamp 1529525674
transform 1 0 20104 0 1 18872
box 0 0 672 896
use LOGIC1_3V  LOGIC1_3V_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 21784 0 -1 20664
box 0 -80 560 976
use BU_3VX2  BU_3VX2_19
timestamp 1529525674
transform 1 0 22344 0 -1 20664
box 0 0 672 896
use BU_3VX2  BU_3VX2_23
timestamp 1529525674
transform 1 0 23016 0 -1 20664
box 0 0 672 896
use BU_3VX2  BU_3VX2_18
timestamp 1529525674
transform 1 0 21560 0 1 18872
box 0 0 672 896
use BU_3VX2  BU_3VX2_21
timestamp 1529525674
transform 1 0 22792 0 1 18872
box 0 0 672 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_4
timestamp 1529525674
transform 1 0 56 0 1 18872
box 0 -80 224 976
use NO2_3VX4  NO2_3VX4_3 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 1400 0 -1 18872
box 0 0 1344 896
use BU_3VX2  BU_3VX2_52
timestamp 1529525674
transform -1 0 2072 0 -1 18872
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_NA3I2_3VX2_1
timestamp 1529525674
transform -1 0 2632 0 -1 18872
box 0 0 560 896
use NA3I2_3VX2  NA3I2_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 3752 0 -1 18872
box 0 0 1120 896
use NA2_3VX0  NA2_3VX0_18
timestamp 1529525674
transform 1 0 3752 0 -1 18872
box 0 0 448 896
use IN_3VX0  IN_3VX0_19
timestamp 1529525674
transform -1 0 4536 0 -1 18872
box 0 0 336 896
use IN_3VX0  IN_3VX0_20
timestamp 1529525674
transform -1 0 4872 0 -1 18872
box 0 0 336 896
use NA3_3VX0  NA3_3VX0_15
timestamp 1529525674
transform -1 0 5432 0 -1 18872
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_16
timestamp 1529525674
transform 1 0 5432 0 -1 18872
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_17
timestamp 1529525674
transform 1 0 5992 0 -1 18872
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_20_0_0
timestamp 1529525674
transform -1 0 7336 0 -1 18872
box 0 0 784 896
use NA3_3VX0  NA3_3VX0_18
timestamp 1529525674
transform -1 0 7896 0 -1 18872
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_13
timestamp 1529525674
transform 1 0 7896 0 -1 18872
box 0 0 3584 896
use BU_3VX2  BU_3VX2_10
timestamp 1529525674
transform 1 0 11480 0 -1 18872
box 0 0 672 896
use BU_3VX2  BU_3VX2_4
timestamp 1529525674
transform -1 0 12824 0 -1 18872
box 0 0 672 896
use BU_3VX2  BU_3VX2_11
timestamp 1529525674
transform -1 0 13496 0 -1 18872
box 0 0 672 896
use MU2_3VX1  MU2_3VX1_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 14728 0 -1 18872
box 0 0 1232 896
use OR2_3VX0  OR2_3VX0_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 14728 0 -1 18872
box 0 0 672 896
use DECAP7_3V  DECAP7_3V_20_1_0
timestamp 1529525674
transform -1 0 16184 0 -1 18872
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_35
timestamp 1529525674
transform -1 0 19768 0 -1 18872
box 0 0 3584 896
use BU_3VX2  BU_3VX2_13
timestamp 1529525674
transform 1 0 19768 0 -1 18872
box 0 0 672 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_10
timestamp 1529525674
transform 1 0 20776 0 1 18872
box 0 -80 224 976
use LOGIC1_3V  LOGIC1_3V_1
timestamp 1529525674
transform 1 0 21000 0 1 18872
box 0 -80 560 976
use LOGIC1_3V  LOGIC1_3V_3
timestamp 1529525674
transform 1 0 22232 0 1 18872
box 0 -80 560 976
use BU_3VX2  BU_3VX2_29
timestamp 1529525674
transform 1 0 20440 0 -1 18872
box 0 0 672 896
use BU_3VX2  BU_3VX2_14
timestamp 1529525674
transform 1 0 21112 0 -1 18872
box 0 0 672 896
use BU_3VX2  BU_3VX2_16
timestamp 1529525674
transform 1 0 21784 0 -1 18872
box 0 0 672 896
use BU_3VX2  BU_3VX2_15
timestamp 1529525674
transform 1 0 22456 0 -1 18872
box 0 0 672 896
use BU_3VX3  BU_3VX3_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 280 0 1 17080
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_NA22_3VX1_3
timestamp 1529525674
transform 1 0 1064 0 1 17080
box 0 0 560 896
use NA22_3VX1  NA22_3VX1_3 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 1624 0 1 17080
box 0 0 784 896
use IN_3VX0  IN_3VX0_18
timestamp 1529525674
transform 1 0 2408 0 1 17080
box 0 0 336 896
use NA2_3VX0  NA2_3VX0_13
timestamp 1529525674
transform 1 0 2744 0 1 17080
box 0 0 448 896
use NA2_3VX0  NA2_3VX0_14
timestamp 1529525674
transform -1 0 3640 0 1 17080
box 0 0 448 896
use NA22_3VX1  NA22_3VX1_4
timestamp 1529525674
transform 1 0 3640 0 1 17080
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_39
timestamp 1529525674
transform 1 0 4424 0 1 17080
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_19_0_0
timestamp 1529525674
transform 1 0 4984 0 1 17080
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_39
timestamp 1529525674
transform 1 0 5768 0 1 17080
box 0 0 3584 896
use OR2_3VX0  OR2_3VX0_2
timestamp 1529525674
transform 1 0 9352 0 1 17080
box 0 0 672 896
use DFRRQ_3VX4  DFRRQ_3VX4_16
timestamp 1529525674
transform 1 0 10024 0 1 17080
box 0 0 3584 896
use DECAP5_3V  DECAP5_3V_1_DFRRQ_3VX4_34
timestamp 1529525674
transform 1 0 13832 0 1 17080
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_34
timestamp 1529525674
transform 1 0 14392 0 1 17080
box 0 0 3584 896
use DECAP7_3V  DECAP7_3V_19_1_0
timestamp 1529525674
transform 1 0 17976 0 1 17080
box 0 0 784 896
use IN_3VX0  IN_3VX0_12
timestamp 1529525674
transform 1 0 18760 0 1 17080
box 0 0 336 896
use LOGIC0_3V  LOGIC0_3V_13
timestamp 1529525674
transform 1 0 19096 0 1 17080
box 0 0 560 896
use DECAP5_3V  DECAP5_3V_0_BU_3VX2_49
timestamp 1529525674
transform 1 0 19656 0 1 17080
box 0 0 560 896
use BU_3VX2  BU_3VX2_49
timestamp 1529525674
transform 1 0 20216 0 1 17080
box 0 0 672 896
use LOGIC0_3V  LOGIC0_3V_4
timestamp 1529525674
transform 1 0 20888 0 1 17080
box 0 0 560 896
use LOGIC1_3V  LOGIC1_3V_4
timestamp 1529525674
transform -1 0 23688 0 -1 18872
box 0 -80 560 976
use BU_3VX2  BU_3VX2_24
timestamp 1529525674
transform 1 0 21448 0 1 17080
box 0 0 672 896
use LOGIC0_3V  LOGIC0_3V_2
timestamp 1529525674
transform 1 0 22120 0 1 17080
box 0 0 560 896
use BU_3VX2  BU_3VX2_20
timestamp 1529525674
transform 1 0 22680 0 1 17080
box 0 0 672 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_1
timestamp 1529525674
transform -1 0 280 0 1 17080
box 0 -80 224 976
use DECAP5_3V  DECAP5_3V_0_IN_3VX4_1
timestamp 1529525674
transform 1 0 56 0 -1 17080
box 0 0 560 896
use IN_3VX4  IN_3VX4_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 616 0 -1 17080
box 0 0 784 896
use NA3_3VX0  NA3_3VX0_13
timestamp 1529525674
transform 1 0 1400 0 -1 17080
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_14
timestamp 1529525674
transform 1 0 1960 0 -1 17080
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_15
timestamp 1529525674
transform 1 0 2520 0 -1 17080
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_NA3_3VX0_12
timestamp 1529525674
transform -1 0 3528 0 -1 17080
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_12
timestamp 1529525674
transform -1 0 4088 0 -1 17080
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_12
timestamp 1529525674
transform -1 0 4536 0 -1 17080
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_1_IN_3VX0_16
timestamp 1529525674
transform -1 0 5320 0 -1 17080
box 0 0 560 896
use IN_3VX0  IN_3VX0_16
timestamp 1529525674
transform -1 0 5656 0 -1 17080
box 0 0 336 896
use NO2_3VX0  NO2_3VX0_10 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 5656 0 -1 17080
box 0 0 448 896
use DECAP7_3V  DECAP7_3V_18_0_0
timestamp 1529525674
transform -1 0 6888 0 -1 17080
box 0 0 784 896
use AO22_3VX1  AO22_3VX1_5 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 7896 0 -1 17080
box 0 0 1008 896
use AO22_3VX1  AO22_3VX1_4
timestamp 1529525674
transform 1 0 7896 0 -1 17080
box 0 0 1008 896
use IN_3VX0  IN_3VX0_15
timestamp 1529525674
transform -1 0 9240 0 -1 17080
box 0 0 336 896
use NA22_3VX1  NA22_3VX1_2
timestamp 1529525674
transform 1 0 9240 0 -1 17080
box 0 0 784 896
use MU2_3VX0  MU2_3VX0_12
timestamp 1529525674
transform 1 0 10024 0 -1 17080
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_DFFRQ_3VX1_9
timestamp 1529525674
transform 1 0 11144 0 -1 17080
box 0 0 560 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_DFRRQ_3VX4_34
timestamp 1529525674
transform 1 0 13608 0 1 17080
box 0 -80 224 976
use DFFRQ_3VX1  DFFRQ_3VX1_9 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 11704 0 -1 17080
box 0 0 3024 896
use MU2_3VX0  MU2_3VX0_5
timestamp 1529525674
transform -1 0 15848 0 -1 17080
box 0 0 1120 896
use MU2_3VX0  MU2_3VX0_6
timestamp 1529525674
transform 1 0 15848 0 -1 17080
box 0 0 1120 896
use DECAP7_3V  DECAP7_3V_18_1_0
timestamp 1529525674
transform 1 0 16968 0 -1 17080
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_DFRSQ_3VX4_5
timestamp 1529525674
transform 1 0 17752 0 -1 17080
box 0 0 560 896
use DFRSQ_3VX4  DFRSQ_3VX4_5
timestamp 1529525674
transform 1 0 18312 0 -1 17080
box 0 0 3360 896
use BU_3VX2  BU_3VX2_27
timestamp 1529525674
transform 1 0 22232 0 -1 17080
box 0 0 672 896
use LOGIC0_3V  LOGIC0_3V_6
timestamp 1529525674
transform 1 0 22904 0 -1 17080
box 0 0 560 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_30
timestamp 1529525674
transform -1 0 616 0 1 15288
box 0 0 560 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_IN_3VX0_16
timestamp 1529525674
transform -1 0 4760 0 -1 17080
box 0 -80 224 976
use DFRRQ_3VX4  DFRRQ_3VX4_30
timestamp 1529525674
transform -1 0 4200 0 1 15288
box 0 0 3584 896
use NA3_3VX2  NA3_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 4200 0 1 15288
box 0 0 1120 896
use NA3_3VX0  NA3_3VX0_11
timestamp 1529525674
transform 1 0 5320 0 1 15288
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_9
timestamp 1529525674
transform 1 0 5880 0 1 15288
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_17_0_0
timestamp 1529525674
transform 1 0 6440 0 1 15288
box 0 0 784 896
use NO2_3VX0  NO2_3VX0_9
timestamp 1529525674
transform 1 0 7224 0 1 15288
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_14
timestamp 1529525674
transform 1 0 7672 0 1 15288
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_14
timestamp 1529525674
transform 1 0 8232 0 1 15288
box 0 0 3584 896
use IN_3VX0  IN_3VX0_13
timestamp 1529525674
transform -1 0 12152 0 1 15288
box 0 0 336 896
use DECAP5_3V  DECAP5_3V_0_MU2_3VX0_26
timestamp 1529525674
transform -1 0 12712 0 1 15288
box 0 0 560 896
use MU2_3VX0  MU2_3VX0_26
timestamp 1529525674
transform -1 0 13832 0 1 15288
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_1_BU_3VX2_1
timestamp 1529525674
transform -1 0 14616 0 1 15288
box 0 0 560 896
use BU_3VX2  BU_3VX2_1
timestamp 1529525674
transform -1 0 15288 0 1 15288
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_DFRSQ_3VX4_4
timestamp 1529525674
transform -1 0 15848 0 1 15288
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_17_1_0
timestamp 1529525674
transform -1 0 16632 0 1 15288
box 0 0 784 896
use DFRSQ_3VX4  DFRSQ_3VX4_4
timestamp 1529525674
transform -1 0 19992 0 1 15288
box 0 0 3360 896
use BU_3VX2  BU_3VX2_22
timestamp 1529525674
transform 1 0 19992 0 1 15288
box 0 0 672 896
use LOGIC0_3V  LOGIC0_3V_10
timestamp 1529525674
transform 1 0 20664 0 1 15288
box 0 0 560 896
use LOGIC1_3V  LOGIC1_3V_5
timestamp 1529525674
transform 1 0 21672 0 -1 17080
box 0 -80 560 976
use BU_3VX2  BU_3VX2_46
timestamp 1529525674
transform 1 0 21224 0 1 15288
box 0 0 672 896
use BU_3VX2  BU_3VX2_45
timestamp 1529525674
transform 1 0 21896 0 1 15288
box 0 0 672 896
use LOGIC0_3V  LOGIC0_3V_8
timestamp 1529525674
transform 1 0 22568 0 1 15288
box 0 0 560 896
use BU_3VX2  BU_3VX2_44
timestamp 1529525674
transform 1 0 23128 0 1 15288
box 0 0 672 896
use BU_3VX2  BU_3VX2_6
timestamp 1529525674
transform 1 0 56 0 -1 15288
box 0 0 672 896
use AO22_3VX1  AO22_3VX1_3
timestamp 1529525674
transform -1 0 1736 0 -1 15288
box 0 0 1008 896
use OA21_3VX2  OA21_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 2968 0 -1 15288
box 0 0 1232 896
use NO2_3VX2  NO2_3VX2_4 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 2968 0 -1 15288
box 0 0 896 896
use NA4_3VX0  NA4_3VX0_6 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 4088 0 -1 15288
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_27
timestamp 1529525674
transform -1 0 5432 0 -1 15288
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_16_0_0
timestamp 1529525674
transform -1 0 6216 0 -1 15288
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_27
timestamp 1529525674
transform -1 0 9800 0 -1 15288
box 0 0 3584 896
use NO22_3VX1  NO22_3VX1_14 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 9800 0 -1 15288
box 0 0 896 896
use DECAP5_3V  DECAP5_3V_0_DFFRQ_3VX1_8
timestamp 1529525674
transform -1 0 11256 0 -1 15288
box 0 0 560 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_BU_3VX2_1
timestamp 1529525674
transform -1 0 14056 0 1 15288
box 0 -80 224 976
use DFFRQ_3VX1  DFFRQ_3VX1_8
timestamp 1529525674
transform -1 0 14280 0 -1 15288
box 0 0 3024 896
use IN_3VX0  IN_3VX0_10
timestamp 1529525674
transform 1 0 14280 0 -1 15288
box 0 0 336 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_3
timestamp 1529525674
transform 1 0 14616 0 -1 15288
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_16_1_0
timestamp 1529525674
transform 1 0 15176 0 -1 15288
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_3
timestamp 1529525674
transform 1 0 15960 0 -1 15288
box 0 0 3584 896
use DECAP5_3V  DECAP5_3V_0_LOGIC0_3V_3
timestamp 1529525674
transform -1 0 20104 0 -1 15288
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_3
timestamp 1529525674
transform -1 0 20664 0 -1 15288
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_5
timestamp 1529525674
transform 1 0 20664 0 -1 15288
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_9
timestamp 1529525674
transform 1 0 21224 0 -1 15288
box 0 0 560 896
use DECAP5_3V  DECAP5_3V_0_BU_3VX2_25
timestamp 1529525674
transform 1 0 21784 0 -1 15288
box 0 0 560 896
use BU_3VX2  BU_3VX2_25
timestamp 1529525674
transform 1 0 22344 0 -1 15288
box 0 0 672 896
use BU_3VX2  BU_3VX2_28
timestamp 1529525674
transform 1 0 23016 0 -1 15288
box 0 0 672 896
use DFFRQ_3VX1  DFFRQ_3VX1_1
timestamp 1529525674
transform 1 0 56 0 1 13496
box 0 0 3024 896
use NO2_3VX0  NO2_3VX0_8
timestamp 1529525674
transform -1 0 3528 0 1 13496
box 0 0 448 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_NA4_3VX0_6
timestamp 1529525674
transform 1 0 3864 0 -1 15288
box 0 -80 224 976
use NO2_3VX2  NO2_3VX2_3
timestamp 1529525674
transform -1 0 4424 0 1 13496
box 0 0 896 896
use NA3_3VX0  NA3_3VX0_21
timestamp 1529525674
transform 1 0 4424 0 1 13496
box 0 0 560 896
use MU2_3VX0  MU2_3VX0_10
timestamp 1529525674
transform 1 0 4984 0 1 13496
box 0 0 1120 896
use IN_3VX0  IN_3VX0_14
timestamp 1529525674
transform -1 0 6440 0 1 13496
box 0 0 336 896
use DECAP7_3V  DECAP7_3V_15_0_0
timestamp 1529525674
transform 1 0 6440 0 1 13496
box 0 0 784 896
use OA22_3VX2  OA22_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 7224 0 1 13496
box 0 0 1344 896
use DECAP5_3V  DECAP5_3V_0_NO3_3VX2_5
timestamp 1529525674
transform -1 0 9128 0 1 13496
box 0 0 560 896
use NO3_3VX2  NO3_3VX2_5 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 10360 0 1 13496
box 0 0 1232 896
use AND2_3VX4  AND2_3VX4_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 10360 0 1 13496
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_BU_3VX3_1
timestamp 1529525674
transform 1 0 11480 0 1 13496
box 0 0 560 896
use BU_3VX3  BU_3VX3_1
timestamp 1529525674
transform 1 0 12040 0 1 13496
box 0 0 784 896
use DFFRQ_3VX1  DFFRQ_3VX1_3
timestamp 1529525674
transform -1 0 15848 0 1 13496
box 0 0 3024 896
use NO22_3VX1  NO22_3VX1_7
timestamp 1529525674
transform -1 0 16744 0 1 13496
box 0 0 896 896
use DECAP7_3V  DECAP7_3V_15_1_0
timestamp 1529525674
transform 1 0 16744 0 1 13496
box 0 0 784 896
use DFRSQ_3VX4  DFRSQ_3VX4_3
timestamp 1529525674
transform 1 0 17752 0 1 13496
box 0 0 3360 896
use DECAP5_3V  DECAP5_3V_0_LOGIC0_3V_12
timestamp 1529525674
transform 1 0 21112 0 1 13496
box 0 0 560 896
use LOGIC0_3V  LOGIC0_3V_12
timestamp 1529525674
transform 1 0 21672 0 1 13496
box 0 0 560 896
use BU_3VX2  BU_3VX2_48
timestamp 1529525674
transform 1 0 22232 0 1 13496
box 0 0 672 896
use LOGIC0_3V  LOGIC0_3V_7
timestamp 1529525674
transform -1 0 23464 0 1 13496
box 0 0 560 896
use BU_3VX2  BU_3VX2_3
timestamp 1529525674
transform 1 0 56 0 -1 13496
box 0 0 672 896
use NO2_3VX2  NO2_3VX2_5
timestamp 1529525674
transform 1 0 728 0 -1 13496
box 0 0 896 896
use NO22_3VX1  NO22_3VX1_15
timestamp 1529525674
transform -1 0 2520 0 -1 13496
box 0 0 896 896
use NA4_3VX2  NA4_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 3976 0 -1 13496
box 0 0 1456 896
use IN_3VX0  IN_3VX0_22
timestamp 1529525674
transform 1 0 3976 0 -1 13496
box 0 0 336 896
use NA2_3VX0  NA2_3VX0_20
timestamp 1529525674
transform 1 0 4312 0 -1 13496
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_29
timestamp 1529525674
transform 1 0 4760 0 -1 13496
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_14_0_0
timestamp 1529525674
transform 1 0 5320 0 -1 13496
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_29
timestamp 1529525674
transform 1 0 6104 0 -1 13496
box 0 0 3584 896
use MU2_3VX0  MU2_3VX0_18
timestamp 1529525674
transform 1 0 9688 0 -1 13496
box 0 0 1120 896
use MU2_3VX0  MU2_3VX0_24
timestamp 1529525674
transform 1 0 10808 0 -1 13496
box 0 0 1120 896
use MU2_3VX0  MU2_3VX0_25
timestamp 1529525674
transform 1 0 11928 0 -1 13496
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_DFFRQ_3VX1_4
timestamp 1529525674
transform -1 0 13608 0 -1 13496
box 0 0 560 896
use DFFRQ_3VX1  DFFRQ_3VX1_4
timestamp 1529525674
transform -1 0 16632 0 -1 13496
box 0 0 3024 896
use DECAP7_3V  DECAP7_3V_14_1_0
timestamp 1529525674
transform 1 0 16632 0 -1 13496
box 0 0 784 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_8
timestamp 1529525674
transform 1 0 17528 0 1 13496
box 0 -80 224 976
use NO3I1_3VX2  NO3I1_3VX2_8 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 17416 0 -1 13496
box 0 0 1456 896
use NO22_3VX1  NO22_3VX1_11
timestamp 1529525674
transform -1 0 19768 0 -1 13496
box 0 0 896 896
use NO22_3VX1  NO22_3VX1_10
timestamp 1529525674
transform 1 0 19992 0 -1 13496
box 0 0 896 896
use NO2I1_3VX1  NO2I1_3VX1_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 20888 0 -1 13496
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_BU_3VX2_41
timestamp 1529525674
transform 1 0 21560 0 -1 13496
box 0 0 560 896
use BU_3VX2  BU_3VX2_41
timestamp 1529525674
transform 1 0 22120 0 -1 13496
box 0 0 672 896
use BU_3VX2  BU_3VX2_42
timestamp 1529525674
transform 1 0 22792 0 -1 13496
box 0 0 672 896
use DFRRQ_3VX4  DFRRQ_3VX4_28
timestamp 1529525674
transform 1 0 56 0 1 11704
box 0 0 3584 896
use MU2_3VX0  MU2_3VX0_11
timestamp 1529525674
transform -1 0 4760 0 1 11704
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_NO3_3VX2_4
timestamp 1529525674
transform 1 0 4760 0 1 11704
box 0 0 560 896
use NO3_3VX2  NO3_3VX2_4
timestamp 1529525674
transform 1 0 5320 0 1 11704
box 0 0 1232 896
use DECAP7_3V  DECAP7_3V_13_0_0
timestamp 1529525674
transform 1 0 6552 0 1 11704
box 0 0 784 896
use NO2_3VX0  NO2_3VX0_13
timestamp 1529525674
transform 1 0 7336 0 1 11704
box 0 0 448 896
use NO2_3VX0  NO2_3VX0_11
timestamp 1529525674
transform -1 0 8232 0 1 11704
box 0 0 448 896
use NO2_3VX0  NO2_3VX0_14
timestamp 1529525674
transform 1 0 8232 0 1 11704
box 0 0 448 896
use NO2_3VX2  NO2_3VX2_6
timestamp 1529525674
transform 1 0 8680 0 1 11704
box 0 0 896 896
use DFFRQ_3VX1  DFFRQ_3VX1_5
timestamp 1529525674
transform -1 0 12600 0 1 11704
box 0 0 3024 896
use MU2_3VX0  MU2_3VX0_17
timestamp 1529525674
transform -1 0 13720 0 1 11704
box 0 0 1120 896
use MU2_3VX0  MU2_3VX0_14
timestamp 1529525674
transform 1 0 13720 0 1 11704
box 0 0 1120 896
use MU2_3VX0  MU2_3VX0_15
timestamp 1529525674
transform 1 0 14840 0 1 11704
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_MU2_3VX0_16
timestamp 1529525674
transform -1 0 16520 0 1 11704
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_13_1_0
timestamp 1529525674
transform -1 0 17304 0 1 11704
box 0 0 784 896
use MU2_3VX0  MU2_3VX0_16
timestamp 1529525674
transform -1 0 18424 0 1 11704
box 0 0 1120 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_NO22_3VX1_10
timestamp 1529525674
transform 1 0 19768 0 -1 13496
box 0 -80 224 976
use NO3I1_3VX2  NO3I1_3VX2_6
timestamp 1529525674
transform 1 0 18424 0 1 11704
box 0 0 1456 896
use NO22_3VX1  NO22_3VX1_9
timestamp 1529525674
transform -1 0 20776 0 1 11704
box 0 0 896 896
use DECAP5_3V  DECAP5_3V_0_NO3I1_3VX2_7
timestamp 1529525674
transform -1 0 21336 0 1 11704
box 0 0 560 896
use NO3I1_3VX2  NO3I1_3VX2_7
timestamp 1529525674
transform -1 0 22792 0 1 11704
box 0 0 1456 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_24
timestamp 1529525674
transform 1 0 56 0 -1 11704
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_24
timestamp 1529525674
transform 1 0 616 0 -1 11704
box 0 0 3584 896
use NO3_3VX0  NO3_3VX0_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 4200 0 -1 11704
box 0 0 672 896
use NO2_3VX0  NO2_3VX0_12
timestamp 1529525674
transform 1 0 4872 0 -1 11704
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_26
timestamp 1529525674
transform -1 0 5880 0 -1 11704
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_12_0_0
timestamp 1529525674
transform -1 0 6664 0 -1 11704
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_26
timestamp 1529525674
transform -1 0 10248 0 -1 11704
box 0 0 3584 896
use DFFRQ_3VX1  DFFRQ_3VX1_7
timestamp 1529525674
transform 1 0 10472 0 -1 11704
box 0 0 3024 896
use MU2_3VX0  MU2_3VX0_22
timestamp 1529525674
transform -1 0 14616 0 -1 11704
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_9
timestamp 1529525674
transform -1 0 15176 0 -1 11704
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_12_1_0
timestamp 1529525674
transform -1 0 15960 0 -1 11704
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_9
timestamp 1529525674
transform -1 0 19544 0 -1 11704
box 0 0 3584 896
use NO3I1_3VX2  NO3I1_3VX2_2
timestamp 1529525674
transform -1 0 21000 0 -1 11704
box 0 0 1456 896
use IN_3VX0  IN_3VX0_11
timestamp 1529525674
transform -1 0 21336 0 -1 11704
box 0 0 336 896
use BU_3VX2  BU_3VX2_40
timestamp 1529525674
transform 1 0 21560 0 -1 11704
box 0 0 672 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_9
timestamp 1529525674
transform 1 0 22792 0 1 11704
box 0 -80 224 976
use LOGIC1_3V  LOGIC1_3V_6
timestamp 1529525674
transform -1 0 23576 0 1 11704
box 0 -80 560 976
use BU_3VX2  BU_3VX2_35
timestamp 1529525674
transform 1 0 22232 0 -1 11704
box 0 0 672 896
use BU_3VX2  BU_3VX2_9
timestamp 1529525674
transform 1 0 56 0 1 9912
box 0 0 672 896
use NA4_3VX0  NA4_3VX0_5
timestamp 1529525674
transform 1 0 952 0 1 9912
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_AND3_3VX2_1
timestamp 1529525674
transform -1 0 2296 0 1 9912
box 0 0 560 896
use AND3_3VX2  AND3_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 3304 0 1 9912
box 0 0 1008 896
use NA2_3VX0  NA2_3VX0_9
timestamp 1529525674
transform -1 0 3752 0 1 9912
box 0 0 448 896
use DFRRQ_3VX4  DFRRQ_3VX4_25
timestamp 1529525674
transform -1 0 7336 0 1 9912
box 0 0 3584 896
use DECAP7_3V  DECAP7_3V_11_0_0
timestamp 1529525674
transform 1 0 7336 0 1 9912
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_DFFRQ_3VX1_6
timestamp 1529525674
transform 1 0 8120 0 1 9912
box 0 0 560 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_DFFRQ_3VX1_7
timestamp 1529525674
transform 1 0 10248 0 -1 11704
box 0 -80 224 976
use DFFRQ_3VX1  DFFRQ_3VX1_6
timestamp 1529525674
transform 1 0 8680 0 1 9912
box 0 0 3024 896
use MU2_3VX0  MU2_3VX0_20
timestamp 1529525674
transform -1 0 12824 0 1 9912
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_MU2_3VX0_21
timestamp 1529525674
transform 1 0 12824 0 1 9912
box 0 0 560 896
use MU2_3VX0  MU2_3VX0_21
timestamp 1529525674
transform 1 0 13384 0 1 9912
box 0 0 1120 896
use AO22_3VX1  AO22_3VX1_1
timestamp 1529525674
transform -1 0 15512 0 1 9912
box 0 0 1008 896
use AO22_3VX1  AO22_3VX1_2
timestamp 1529525674
transform -1 0 16520 0 1 9912
box 0 0 1008 896
use DECAP7_3V  DECAP7_3V_11_1_0
timestamp 1529525674
transform -1 0 17304 0 1 9912
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_NO3I2_3VX1_3
timestamp 1529525674
transform -1 0 17864 0 1 9912
box 0 0 560 896
use NO3I2_3VX1  NO3I2_3VX1_3 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 18648 0 1 9912
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_NO22_3VX1_5
timestamp 1529525674
transform 1 0 18648 0 1 9912
box 0 0 560 896
use NO22_3VX1  NO22_3VX1_5
timestamp 1529525674
transform 1 0 19208 0 1 9912
box 0 0 896 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_BU_3VX2_40
timestamp 1529525674
transform 1 0 21336 0 -1 11704
box 0 -80 224 976
use LOGIC1_3V  LOGIC1_3V_7
timestamp 1529525674
transform 1 0 22904 0 -1 11704
box 0 -80 560 976
use DFRRQ_3VX4  DFRRQ_3VX4_1
timestamp 1529525674
transform -1 0 23688 0 1 9912
box 0 0 3584 896
use NA2I1_3VX1  NA2I1_3VX1_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 56 0 -1 9912
box 0 0 672 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_2
timestamp 1529525674
transform 1 0 728 0 1 9912
box 0 -80 224 976
use NA22_3VX1  NA22_3VX1_10
timestamp 1529525674
transform 1 0 728 0 -1 9912
box 0 0 784 896
use NO3I2_3VX1  NO3I2_3VX1_4
timestamp 1529525674
transform -1 0 2296 0 -1 9912
box 0 0 784 896
use IN_3VX0  IN_3VX0_26
timestamp 1529525674
transform -1 0 2632 0 -1 9912
box 0 0 336 896
use ON31_3VX2  ON31_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 4088 0 -1 9912
box 0 0 1456 896
use NA2I1_3VX1  NA2I1_3VX1_1
timestamp 1529525674
transform -1 0 4760 0 -1 9912
box 0 0 672 896
use DECAP7_3V  DECAP7_3V_10_0_0
timestamp 1529525674
transform 1 0 4760 0 -1 9912
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_19
timestamp 1529525674
transform 1 0 5544 0 -1 9912
box 0 0 3584 896
use BU_3VX2  BU_3VX2_2
timestamp 1529525674
transform 1 0 9128 0 -1 9912
box 0 0 672 896
use BU_3VX2  BU_3VX2_8
timestamp 1529525674
transform -1 0 10696 0 -1 9912
box 0 0 672 896
use MU2_3VX0  MU2_3VX0_19
timestamp 1529525674
transform 1 0 10696 0 -1 9912
box 0 0 1120 896
use MU2_3VX0  MU2_3VX0_23
timestamp 1529525674
transform -1 0 12936 0 -1 9912
box 0 0 1120 896
use AN22_3VX2  AN22_3VX2_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 14392 0 -1 9912
box 0 0 1456 896
use NA3_3VX0  NA3_3VX0_3
timestamp 1529525674
transform 1 0 14392 0 -1 9912
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_6
timestamp 1529525674
transform -1 0 15400 0 -1 9912
box 0 0 448 896
use NO22_3VX1  NO22_3VX1_4
timestamp 1529525674
transform 1 0 15400 0 -1 9912
box 0 0 896 896
use DECAP7_3V  DECAP7_3V_10_1_0
timestamp 1529525674
transform 1 0 16296 0 -1 9912
box 0 0 784 896
use NO22_3VX1  NO22_3VX1_3
timestamp 1529525674
transform 1 0 17080 0 -1 9912
box 0 0 896 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_8
timestamp 1529525674
transform -1 0 18536 0 -1 9912
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_8
timestamp 1529525674
transform -1 0 22120 0 -1 9912
box 0 0 3584 896
use BU_3VX2  BU_3VX2_47
timestamp 1529525674
transform 1 0 22120 0 -1 9912
box 0 0 672 896
use BU_3VX2  BU_3VX2_43
timestamp 1529525674
transform 1 0 22792 0 -1 9912
box 0 0 672 896
use MU2_3VX1  MU2_3VX1_5
timestamp 1529525674
transform -1 0 1288 0 1 8120
box 0 0 1232 896
use DECAP5_3V  DECAP5_3V_0_OA22_3VX2_2
timestamp 1529525674
transform -1 0 1848 0 1 8120
box 0 0 560 896
use OA22_3VX2  OA22_3VX2_2
timestamp 1529525674
transform -1 0 3192 0 1 8120
box 0 0 1344 896
use IN_3VX0  IN_3VX0_25
timestamp 1529525674
transform -1 0 3528 0 1 8120
box 0 0 336 896
use NA3_3VX0  NA3_3VX0_10
timestamp 1529525674
transform -1 0 4088 0 1 8120
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_11
timestamp 1529525674
transform -1 0 4536 0 1 8120
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_NA2_3VX0_29
timestamp 1529525674
transform 1 0 4536 0 1 8120
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_29
timestamp 1529525674
transform 1 0 5096 0 1 8120
box 0 0 448 896
use NA3_3VX0  NA3_3VX0_24
timestamp 1529525674
transform -1 0 6104 0 1 8120
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_9_0_0
timestamp 1529525674
transform 1 0 6104 0 1 8120
box 0 0 784 896
use NA2_3VX0  NA2_3VX0_10
timestamp 1529525674
transform 1 0 6888 0 1 8120
box 0 0 448 896
use NA2_3VX0  NA2_3VX0_23
timestamp 1529525674
transform -1 0 7784 0 1 8120
box 0 0 448 896
use NO2_3VX4  NO2_3VX4_2
timestamp 1529525674
transform 1 0 7784 0 1 8120
box 0 0 1344 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_3
timestamp 1529525674
transform -1 0 10024 0 -1 9912
box 0 -80 224 976
use NO2_3VX2  NO2_3VX2_2
timestamp 1529525674
transform 1 0 9128 0 1 8120
box 0 0 896 896
use DFRRQ_3VX4  DFRRQ_3VX4_7
timestamp 1529525674
transform 1 0 10024 0 1 8120
box 0 0 3584 896
use AN22_3VX2  AN22_3VX2_1
timestamp 1529525674
transform -1 0 15064 0 1 8120
box 0 0 1456 896
use IN_3VX0  IN_3VX0_9
timestamp 1529525674
transform 1 0 15064 0 1 8120
box 0 0 336 896
use NA3_3VX0  NA3_3VX0_2
timestamp 1529525674
transform -1 0 15960 0 1 8120
box 0 0 560 896
use NO2_3VX0  NO2_3VX0_3
timestamp 1529525674
transform 1 0 15960 0 1 8120
box 0 0 448 896
use DECAP7_3V  DECAP7_3V_9_1_0
timestamp 1529525674
transform -1 0 17192 0 1 8120
box 0 0 784 896
use NO2_3VX0  NO2_3VX0_5
timestamp 1529525674
transform -1 0 17640 0 1 8120
box 0 0 448 896
use NO22_3VX1  NO22_3VX1_2
timestamp 1529525674
transform -1 0 18536 0 1 8120
box 0 0 896 896
use BU_3VX2  BU_3VX2_55
timestamp 1529525674
transform 1 0 18536 0 1 8120
box 0 0 672 896
use NO2_3VX0  NO2_3VX0_4
timestamp 1529525674
transform -1 0 19656 0 1 8120
box 0 0 448 896
use BU_3VX2  BU_3VX2_5
timestamp 1529525674
transform 1 0 19656 0 1 8120
box 0 0 672 896
use NO2I1_3VX4  NO2I1_3VX4_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 20328 0 1 8120
box 0 0 1568 896
use LOGIC0_3V  LOGIC0_3V_11
timestamp 1529525674
transform 1 0 21896 0 1 8120
box 0 0 560 896
use DECAP5_3V  DECAP5_3V_0_BU_3VX2_57
timestamp 1529525674
transform 1 0 22456 0 1 8120
box 0 0 560 896
use BU_3VX2  BU_3VX2_57
timestamp 1529525674
transform 1 0 23016 0 1 8120
box 0 0 672 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_DFRRQ_3VX4_12
timestamp 1529525674
transform 1 0 56 0 -1 8120
box 0 -80 224 976
use DECAP5_3V  DECAP5_3V_1_DFRRQ_3VX4_12
timestamp 1529525674
transform 1 0 280 0 -1 8120
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_12
timestamp 1529525674
transform 1 0 840 0 -1 8120
box 0 0 3584 896
use AO31_3VX1  AO31_3VX1_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 4424 0 -1 8120
box 0 0 1120 896
use NA3_3VX0  NA3_3VX0_23
timestamp 1529525674
transform -1 0 6104 0 -1 8120
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_8_0_0
timestamp 1529525674
transform -1 0 6888 0 -1 8120
box 0 0 784 896
use NA4_3VX2  NA4_3VX2_2
timestamp 1529525674
transform -1 0 8344 0 -1 8120
box 0 0 1456 896
use BU_3VX3  BU_3VX3_3
timestamp 1529525674
transform -1 0 9128 0 -1 8120
box 0 0 784 896
use IN_3VX1  IN_3VX1_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 9128 0 -1 8120
box 0 0 336 896
use BU_3VX2  BU_3VX2_7
timestamp 1529525674
transform 1 0 9464 0 -1 8120
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_DFFRQ_3VX1_2
timestamp 1529525674
transform 1 0 10136 0 -1 8120
box 0 0 560 896
use DFFRQ_3VX1  DFFRQ_3VX1_2
timestamp 1529525674
transform 1 0 10696 0 -1 8120
box 0 0 3024 896
use DECAP5_3V  DECAP5_3V_0_NA22_3VX1_1
timestamp 1529525674
transform -1 0 14280 0 -1 8120
box 0 0 560 896
use NA22_3VX1  NA22_3VX1_1
timestamp 1529525674
transform -1 0 15064 0 -1 8120
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_NA3_3VX0_4
timestamp 1529525674
transform -1 0 15624 0 -1 8120
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_4
timestamp 1529525674
transform -1 0 16184 0 -1 8120
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_7
timestamp 1529525674
transform -1 0 16632 0 -1 8120
box 0 0 448 896
use DECAP7_3V  DECAP7_3V_8_1_0
timestamp 1529525674
transform -1 0 17416 0 -1 8120
box 0 0 784 896
use NA3_3VX0  NA3_3VX0_1
timestamp 1529525674
transform -1 0 17976 0 -1 8120
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_5
timestamp 1529525674
transform -1 0 18536 0 -1 8120
box 0 0 560 896
use DECAP5_3V  DECAP5_3V_0_NO2_3VX0_2
timestamp 1529525674
transform -1 0 19096 0 -1 8120
box 0 0 560 896
use NO2_3VX0  NO2_3VX0_2
timestamp 1529525674
transform -1 0 19544 0 -1 8120
box 0 0 448 896
use NA2_3VX4  NA2_3VX4_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 21000 0 -1 8120
box 0 0 1456 896
use NO22_3VX1  NO22_3VX1_6
timestamp 1529525674
transform 1 0 21224 0 -1 8120
box 0 0 896 896
use NO3I1_3VX2  NO3I1_3VX2_3
timestamp 1529525674
transform -1 0 23576 0 -1 8120
box 0 0 1456 896
use DECAP5_3V  DECAP5_3V_1_DFRRQ_3VX4_23
timestamp 1529525674
transform 1 0 280 0 1 6328
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_23
timestamp 1529525674
transform 1 0 840 0 1 6328
box 0 0 3584 896
use NA22_3VX1  NA22_3VX1_6
timestamp 1529525674
transform -1 0 5208 0 1 6328
box 0 0 784 896
use OA31_3VX1  OA31_3VX1_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 6216 0 1 6328
box 0 0 1008 896
use DECAP7_3V  DECAP7_3V_7_0_0
timestamp 1529525674
transform -1 0 7000 0 1 6328
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_NA22_3VX1_5
timestamp 1529525674
transform -1 0 7560 0 1 6328
box 0 0 560 896
use NA22_3VX1  NA22_3VX1_5
timestamp 1529525674
transform -1 0 8344 0 1 6328
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_22
timestamp 1529525674
transform -1 0 11928 0 1 6328
box 0 0 3584 896
use NA2I1_3VX1  NA2I1_3VX1_3
timestamp 1529525674
transform 1 0 11928 0 1 6328
box 0 0 672 896
use NA2_3VX0  NA2_3VX0_36
timestamp 1529525674
transform -1 0 13048 0 1 6328
box 0 0 448 896
use MU2_3VX0  MU2_3VX0_13
timestamp 1529525674
transform 1 0 13048 0 1 6328
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_NA3_3VX0_25
timestamp 1529525674
transform -1 0 14728 0 1 6328
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_25
timestamp 1529525674
transform -1 0 15288 0 1 6328
box 0 0 560 896
use NA4_3VX0  NA4_3VX0_2
timestamp 1529525674
transform 1 0 15512 0 1 6328
box 0 0 784 896
use NA2_3VX0  NA2_3VX0_5
timestamp 1529525674
transform -1 0 16744 0 1 6328
box 0 0 448 896
use DECAP7_3V  DECAP7_3V_7_1_0
timestamp 1529525674
transform 1 0 16744 0 1 6328
box 0 0 784 896
use IN_3VX1  IN_3VX1_1
timestamp 1529525674
transform 1 0 17528 0 1 6328
box 0 0 336 896
use NA2_3VX0  NA2_3VX0_4
timestamp 1529525674
transform -1 0 18312 0 1 6328
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_NO2_3VX0_6
timestamp 1529525674
transform 1 0 18312 0 1 6328
box 0 0 560 896
use NO2_3VX0  NO2_3VX0_6
timestamp 1529525674
transform 1 0 18872 0 1 6328
box 0 0 448 896
use NA2_3VX0  NA2_3VX0_8
timestamp 1529525674
transform -1 0 19768 0 1 6328
box 0 0 448 896
use NO22_3VX1  NO22_3VX1_8
timestamp 1529525674
transform -1 0 20664 0 1 6328
box 0 0 896 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_6
timestamp 1529525674
transform -1 0 21224 0 -1 8120
box 0 -80 224 976
use AND2_3VX0  AND2_3VX0_1
timestamp 1529525674
transform 1 0 20664 0 1 6328
box 0 0 672 896
use NO22_3VX1  NO22_3VX1_12
timestamp 1529525674
transform 1 0 21336 0 1 6328
box 0 0 896 896
use DECAP5_3V  DECAP5_3V_0_BU_3VX2_33
timestamp 1529525674
transform 1 0 22232 0 1 6328
box 0 0 560 896
use BU_3VX2  BU_3VX2_33
timestamp 1529525674
transform 1 0 22792 0 1 6328
box 0 0 672 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_DFRRQ_3VX4_23
timestamp 1529525674
transform 1 0 56 0 1 6328
box 0 -80 224 976
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_20
timestamp 1529525674
transform 1 0 56 0 -1 6328
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_20
timestamp 1529525674
transform 1 0 616 0 -1 6328
box 0 0 3584 896
use IN_3VX0  IN_3VX0_24
timestamp 1529525674
transform -1 0 4536 0 -1 6328
box 0 0 336 896
use NA22_3VX1  NA22_3VX1_8
timestamp 1529525674
transform 1 0 4536 0 -1 6328
box 0 0 784 896
use NA22_3VX1  NA22_3VX1_9
timestamp 1529525674
transform 1 0 5320 0 -1 6328
box 0 0 784 896
use DECAP7_3V  DECAP7_3V_6_0_0
timestamp 1529525674
transform -1 0 6888 0 -1 6328
box 0 0 784 896
use NA2_3VX0  NA2_3VX0_30
timestamp 1529525674
transform -1 0 7336 0 -1 6328
box 0 0 448 896
use NA2_3VX2  NA2_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 8120 0 -1 6328
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_38
timestamp 1529525674
transform 1 0 8120 0 -1 6328
box 0 0 3584 896
use DECAP5_3V  DECAP5_3V_0_NA3_3VX0_8
timestamp 1529525674
transform 1 0 11704 0 -1 6328
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_8
timestamp 1529525674
transform 1 0 12264 0 -1 6328
box 0 0 560 896
use NO3I1_3VX2  NO3I1_3VX2_4
timestamp 1529525674
transform 1 0 12824 0 -1 6328
box 0 0 1456 896
use NA2_3VX0  NA2_3VX0_3
timestamp 1529525674
transform 1 0 14280 0 -1 6328
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_NO3I1_3VX2_5
timestamp 1529525674
transform 1 0 14728 0 -1 6328
box 0 0 560 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_NA4_3VX0_2
timestamp 1529525674
transform 1 0 15288 0 1 6328
box 0 -80 224 976
use NO3I1_3VX2  NO3I1_3VX2_5
timestamp 1529525674
transform 1 0 15288 0 -1 6328
box 0 0 1456 896
use DECAP7_3V  DECAP7_3V_6_1_0
timestamp 1529525674
transform 1 0 16744 0 -1 6328
box 0 0 784 896
use BU_3VX2  BU_3VX2_54
timestamp 1529525674
transform 1 0 17528 0 -1 6328
box 0 0 672 896
use NO2_3VX0  NO2_3VX0_7
timestamp 1529525674
transform 1 0 18200 0 -1 6328
box 0 0 448 896
use NO22_3VX1  NO22_3VX1_13
timestamp 1529525674
transform -1 0 19544 0 -1 6328
box 0 0 896 896
use DECAP5_3V  DECAP5_3V_0_DFRSQ_3VX4_2
timestamp 1529525674
transform -1 0 20104 0 -1 6328
box 0 0 560 896
use DFRSQ_3VX4  DFRSQ_3VX4_2
timestamp 1529525674
transform -1 0 23464 0 -1 6328
box 0 0 3360 896
use NA2_3VX0  NA2_3VX0_34
timestamp 1529525674
transform -1 0 504 0 1 4536
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_AO31_3VX1_4
timestamp 1529525674
transform -1 0 1064 0 1 4536
box 0 0 560 896
use AO31_3VX1  AO31_3VX1_4
timestamp 1529525674
transform -1 0 2184 0 1 4536
box 0 0 1120 896
use NA4_3VX0  NA4_3VX0_4
timestamp 1529525674
transform -1 0 2968 0 1 4536
box 0 0 784 896
use NA2_3VX0  NA2_3VX0_25
timestamp 1529525674
transform -1 0 3416 0 1 4536
box 0 0 448 896
use IN_3VX0  IN_3VX0_23
timestamp 1529525674
transform 1 0 3416 0 1 4536
box 0 0 336 896
use OA31_3VX1  OA31_3VX1_2
timestamp 1529525674
transform 1 0 4200 0 1 4536
box 0 0 1008 896
use NA2_3VX0  NA2_3VX0_26
timestamp 1529525674
transform 1 0 5208 0 1 4536
box 0 0 448 896
use NA4_3VX0  NA4_3VX0_3
timestamp 1529525674
transform 1 0 5656 0 1 4536
box 0 0 784 896
use DECAP7_3V  DECAP7_3V_5_0_0
timestamp 1529525674
transform 1 0 6440 0 1 4536
box 0 0 784 896
use NA2_3VX0  NA2_3VX0_27
timestamp 1529525674
transform 1 0 7224 0 1 4536
box 0 0 448 896
use AO31_3VX1  AO31_3VX1_1
timestamp 1529525674
transform -1 0 8792 0 1 4536
box 0 0 1120 896
use MU2_3VX0  MU2_3VX0_8
timestamp 1529525674
transform -1 0 9912 0 1 4536
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_MU2_3VX0_9
timestamp 1529525674
transform -1 0 10472 0 1 4536
box 0 0 560 896
use MU2_3VX0  MU2_3VX0_9
timestamp 1529525674
transform -1 0 11592 0 1 4536
box 0 0 1120 896
use MU2_3VX0  MU2_3VX0_3
timestamp 1529525674
transform -1 0 12712 0 1 4536
box 0 0 1120 896
use IN_3VX0  IN_3VX0_6
timestamp 1529525674
transform -1 0 13048 0 1 4536
box 0 0 336 896
use NO3_3VX2  NO3_3VX2_3
timestamp 1529525674
transform 1 0 13048 0 1 4536
box 0 0 1232 896
use NO2_3VX2  NO2_3VX2_1
timestamp 1529525674
transform -1 0 15176 0 1 4536
box 0 0 896 896
use NO3_3VX2  NO3_3VX2_2
timestamp 1529525674
transform -1 0 16408 0 1 4536
box 0 0 1232 896
use DECAP7_3V  DECAP7_3V_5_1_0
timestamp 1529525674
transform 1 0 16408 0 1 4536
box 0 0 784 896
use AND2_3VX1  AND2_3VX1_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 17192 0 1 4536
box 0 0 672 896
use NO22_3VX1  NO22_3VX1_1
timestamp 1529525674
transform 1 0 17864 0 1 4536
box 0 0 896 896
use IN_3VX0  IN_3VX0_8
timestamp 1529525674
transform -1 0 19096 0 1 4536
box 0 0 336 896
use DFRRQ_3VX4  DFRRQ_3VX4_4
timestamp 1529525674
transform 1 0 19320 0 1 4536
box 0 0 3584 896
use BU_3VX2  BU_3VX2_34
timestamp 1529525674
transform 1 0 22904 0 1 4536
box 0 0 672 896
use AO21_3VX1  AO21_3VX1_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 56 0 -1 4536
box 0 0 896 896
use AO22_3VX1  AO22_3VX1_8
timestamp 1529525674
transform -1 0 1960 0 -1 4536
box 0 0 1008 896
use NA2_3VX0  NA2_3VX0_31
timestamp 1529525674
transform 1 0 1960 0 -1 4536
box 0 0 448 896
use NA22_3VX1  NA22_3VX1_7
timestamp 1529525674
transform -1 0 3192 0 -1 4536
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_NA2_3VX0_32
timestamp 1529525674
transform 1 0 3192 0 -1 4536
box 0 0 560 896
use IN_3VX2  IN_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 3752 0 1 4536
box 0 -80 448 976
use NA2_3VX0  NA2_3VX0_32
timestamp 1529525674
transform 1 0 3752 0 -1 4536
box 0 0 448 896
use IN_3VX0  IN_3VX0_17
timestamp 1529525674
transform 1 0 4200 0 -1 4536
box 0 0 336 896
use NA2_3VX0  NA2_3VX0_28
timestamp 1529525674
transform 1 0 4536 0 -1 4536
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_37
timestamp 1529525674
transform 1 0 4984 0 -1 4536
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_4_0_0
timestamp 1529525674
transform 1 0 5544 0 -1 4536
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_37
timestamp 1529525674
transform 1 0 6328 0 -1 4536
box 0 0 3584 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_5
timestamp 1529525674
transform 1 0 9912 0 -1 4536
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_5
timestamp 1529525674
transform 1 0 10472 0 -1 4536
box 0 0 3584 896
use NO3I2_3VX1  NO3I2_3VX1_2
timestamp 1529525674
transform 1 0 14056 0 -1 4536
box 0 0 784 896
use OR2_3VX1  OR2_3VX1_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 14840 0 -1 4536
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_NO3_3VX2_1
timestamp 1529525674
transform 1 0 15512 0 -1 4536
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_4_1_0
timestamp 1529525674
transform 1 0 16072 0 -1 4536
box 0 0 784 896
use NO3_3VX2  NO3_3VX2_1
timestamp 1529525674
transform 1 0 16856 0 -1 4536
box 0 0 1232 896
use NA3I2_3VX1  NA3I2_3VX1_3
timestamp 1529525674
transform -1 0 18872 0 -1 4536
box 0 0 784 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_DFRRQ_3VX4_4
timestamp 1529525674
transform 1 0 19096 0 1 4536
box 0 -80 224 976
use DFRSQ_3VX4  DFRSQ_3VX4_1
timestamp 1529525674
transform 1 0 18872 0 -1 4536
box 0 0 3360 896
use BU_3VX2  BU_3VX2_50
timestamp 1529525674
transform 1 0 22232 0 -1 4536
box 0 0 672 896
use BU_3VX2  BU_3VX2_26
timestamp 1529525674
transform 1 0 22904 0 -1 4536
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_MU2_3VX1_4
timestamp 1529525674
transform -1 0 616 0 1 2744
box 0 0 560 896
use MU2_3VX1  MU2_3VX1_4
timestamp 1529525674
transform -1 0 1848 0 1 2744
box 0 0 1232 896
use AO22_3VX1  AO22_3VX1_7
timestamp 1529525674
transform -1 0 2856 0 1 2744
box 0 0 1008 896
use DECAP5_3V  DECAP5_3V_0_AO31_3VX1_3
timestamp 1529525674
transform -1 0 3416 0 1 2744
box 0 0 560 896
use AO31_3VX1  AO31_3VX1_3
timestamp 1529525674
transform -1 0 4536 0 1 2744
box 0 0 1120 896
use NA4_3VX2  NA4_3VX2_3
timestamp 1529525674
transform -1 0 5992 0 1 2744
box 0 0 1456 896
use DECAP5_3V  DECAP5_3V_0_NA2_3VX0_24
timestamp 1529525674
transform 1 0 5992 0 1 2744
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_3_0_0
timestamp 1529525674
transform 1 0 6552 0 1 2744
box 0 0 784 896
use NA2_3VX0  NA2_3VX0_24
timestamp 1529525674
transform 1 0 7336 0 1 2744
box 0 0 448 896
use NA3_3VX0  NA3_3VX0_22
timestamp 1529525674
transform 1 0 7784 0 1 2744
box 0 0 560 896
use NO2_3VX0  NO2_3VX0_15
timestamp 1529525674
transform -1 0 9016 0 1 2744
box 0 0 448 896
use DFRRQ_3VX4  DFRRQ_3VX4_11
timestamp 1529525674
transform 1 0 9016 0 1 2744
box 0 0 3584 896
use MU2_3VX0  MU2_3VX0_1
timestamp 1529525674
transform -1 0 13720 0 1 2744
box 0 0 1120 896
use NA2I1_3VX2  NA2I1_3VX2_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 14728 0 1 2744
box 0 0 1008 896
use NA2I1_3VX2  NA2I1_3VX2_3
timestamp 1529525674
transform 1 0 14728 0 1 2744
box 0 0 1008 896
use NA2_3VX0  NA2_3VX0_2
timestamp 1529525674
transform 1 0 15736 0 1 2744
box 0 0 448 896
use DECAP7_3V  DECAP7_3V_3_1_0
timestamp 1529525674
transform 1 0 16184 0 1 2744
box 0 0 784 896
use OR4_3VX1  OR4_3VX1_4 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 16968 0 1 2744
box 0 0 1232 896
use OR4_3VX1  OR4_3VX1_3
timestamp 1529525674
transform 1 0 18200 0 1 2744
box 0 0 1232 896
use DECAP5_3V  DECAP5_3V_0_OR4_3VX1_1
timestamp 1529525674
transform 1 0 19432 0 1 2744
box 0 0 560 896
use OR4_3VX1  OR4_3VX1_1
timestamp 1529525674
transform 1 0 19992 0 1 2744
box 0 0 1232 896
use IN_3VX0  IN_3VX0_2
timestamp 1529525674
transform -1 0 21560 0 1 2744
box 0 0 336 896
use IN_3VX0  IN_3VX0_4
timestamp 1529525674
transform -1 0 21896 0 1 2744
box 0 0 336 896
use BU_3VX2  BU_3VX2_39
timestamp 1529525674
transform -1 0 22568 0 1 2744
box 0 0 672 896
use BU_3VX2  BU_3VX2_51
timestamp 1529525674
transform 1 0 22568 0 1 2744
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_21
timestamp 1529525674
transform 1 0 56 0 -1 2744
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_21
timestamp 1529525674
transform 1 0 616 0 -1 2744
box 0 0 3584 896
use NA3I2_3VX1  NA3I2_3VX1_5
timestamp 1529525674
transform -1 0 4984 0 -1 2744
box 0 0 784 896
use NO3I1_3VX2  NO3I1_3VX2_9
timestamp 1529525674
transform -1 0 6440 0 -1 2744
box 0 0 1456 896
use DECAP7_3V  DECAP7_3V_2_0_0
timestamp 1529525674
transform -1 0 7224 0 -1 2744
box 0 0 784 896
use NO2I1_3VX2  NO2I1_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 8232 0 -1 2744
box 0 0 1008 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_0_NO2_3VX0_15
timestamp 1529525674
transform -1 0 8568 0 1 2744
box 0 -80 224 976
use AO22_3VX1  AO22_3VX1_6
timestamp 1529525674
transform -1 0 9240 0 -1 2744
box 0 0 1008 896
use NA2_3VX0  NA2_3VX0_22
timestamp 1529525674
transform -1 0 9688 0 -1 2744
box 0 0 448 896
use NA22_3VX1  NA22_3VX1_11
timestamp 1529525674
transform 1 0 9688 0 -1 2744
box 0 0 784 896
use NA2_3VX0  NA2_3VX0_21
timestamp 1529525674
transform -1 0 10920 0 -1 2744
box 0 0 448 896
use MU2_3VX4  MU2_3VX4_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 10920 0 -1 2744
box 0 0 1680 896
use DECAP5_3V  DECAP5_3V_0_NO2_3VX0_1
timestamp 1529525674
transform 1 0 12600 0 -1 2744
box 0 0 560 896
use NO2_3VX0  NO2_3VX0_1
timestamp 1529525674
transform 1 0 13160 0 -1 2744
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_NA2_3VX0_1
timestamp 1529525674
transform -1 0 14168 0 -1 2744
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_1
timestamp 1529525674
transform -1 0 14616 0 -1 2744
box 0 0 448 896
use IN_3VX0  IN_3VX0_7
timestamp 1529525674
transform 1 0 14616 0 -1 2744
box 0 0 336 896
use NA3I2_3VX1  NA3I2_3VX1_2
timestamp 1529525674
transform 1 0 14952 0 -1 2744
box 0 0 784 896
use NA3_3VX0  NA3_3VX0_6
timestamp 1529525674
transform 1 0 15736 0 -1 2744
box 0 0 560 896
use NA3_3VX0  NA3_3VX0_7
timestamp 1529525674
transform 1 0 16296 0 -1 2744
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_2_1_0
timestamp 1529525674
transform 1 0 16856 0 -1 2744
box 0 0 784 896
use NA4_3VX0  NA4_3VX0_1
timestamp 1529525674
transform 1 0 17640 0 -1 2744
box 0 0 784 896
use IN_3VX0  IN_3VX0_1
timestamp 1529525674
transform 1 0 18424 0 -1 2744
box 0 0 336 896
use BU_3VX2  BU_3VX2_36
timestamp 1529525674
transform 1 0 18760 0 -1 2744
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_6
timestamp 1529525674
transform -1 0 19992 0 -1 2744
box 0 0 560 896
use ANTENNACELLNP2_3V  ANTENNACELLNP2_3V_5
timestamp 1529525674
transform -1 0 23464 0 1 2744
box 0 -80 224 976
use DFRRQ_3VX4  DFRRQ_3VX4_6
timestamp 1529525674
transform -1 0 23576 0 -1 2744
box 0 0 3584 896
use OR4_3VX2  OR4_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 56 0 1 952
box 0 0 1456 896
use MU2_3VX1  MU2_3VX1_3
timestamp 1529525674
transform -1 0 2744 0 1 952
box 0 0 1232 896
use MU2_3VX1  MU2_3VX1_2
timestamp 1529525674
transform -1 0 3976 0 1 952
box 0 0 1232 896
use NA2_3VX0  NA2_3VX0_33
timestamp 1529525674
transform 1 0 3976 0 1 952
box 0 0 448 896
use DECAP5_3V  DECAP5_3V_0_NA2_3VX0_35
timestamp 1529525674
transform 1 0 4424 0 1 952
box 0 0 560 896
use NA2_3VX0  NA2_3VX0_35
timestamp 1529525674
transform 1 0 4984 0 1 952
box 0 0 448 896
use NA3_3VX2  NA3_3VX2_2
timestamp 1529525674
transform 1 0 5432 0 1 952
box 0 0 1120 896
use DECAP7_3V  DECAP7_3V_1_0_0
timestamp 1529525674
transform 1 0 6552 0 1 952
box 0 0 784 896
use MU2_3VX4  MU2_3VX4_3
timestamp 1529525674
transform 1 0 7336 0 1 952
box 0 0 1680 896
use DECAP5_3V  DECAP5_3V_0_MU2_3VX4_2
timestamp 1529525674
transform 1 0 9016 0 1 952
box 0 0 560 896
use MU2_3VX4  MU2_3VX4_2
timestamp 1529525674
transform 1 0 9576 0 1 952
box 0 0 1680 896
use NO3I1_3VX2  NO3I1_3VX2_1
timestamp 1529525674
transform 1 0 11256 0 1 952
box 0 0 1456 896
use OR2_3VX1  OR2_3VX1_2
timestamp 1529525674
transform 1 0 12712 0 1 952
box 0 0 672 896
use OR2_3VX2  OR2_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform 1 0 13384 0 1 952
box 0 0 896 896
use NA3I2_3VX1  NA3I2_3VX1_1
timestamp 1529525674
transform -1 0 15064 0 1 952
box 0 0 784 896
use IN_3VX0  IN_3VX0_5
timestamp 1529525674
transform 1 0 15064 0 1 952
box 0 0 336 896
use DECAP5_3V  DECAP5_3V_0_NO3I2_3VX1_1
timestamp 1529525674
transform 1 0 15400 0 1 952
box 0 0 560 896
use NO3I2_3VX1  NO3I2_3VX1_1
timestamp 1529525674
transform 1 0 15960 0 1 952
box 0 0 784 896
use DECAP7_3V  DECAP7_3V_1_1_0
timestamp 1529525674
transform 1 0 16744 0 1 952
box 0 0 784 896
use MU2_3VX0  MU2_3VX0_2
timestamp 1529525674
transform 1 0 17528 0 1 952
box 0 0 1120 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_10
timestamp 1529525674
transform 1 0 18648 0 1 952
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_10
timestamp 1529525674
transform 1 0 19208 0 1 952
box 0 0 3584 896
use BU_3VX2  BU_3VX2_12
timestamp 1529525674
transform 1 0 22792 0 1 952
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_17
timestamp 1529525674
transform 1 0 56 0 -1 952
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_17
timestamp 1529525674
transform 1 0 616 0 -1 952
box 0 0 3584 896
use AND2_3VX2  AND2_3VX2_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/D_CELLS_3V
timestamp 1529525674
transform -1 0 4984 0 -1 952
box 0 0 784 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_18
timestamp 1529525674
transform 1 0 4984 0 -1 952
box 0 0 560 896
use DECAP7_3V  DECAP7_3V_0_0_0
timestamp 1529525674
transform 1 0 5544 0 -1 952
box 0 0 784 896
use DFRRQ_3VX4  DFRRQ_3VX4_18
timestamp 1529525674
transform 1 0 6328 0 -1 952
box 0 0 3584 896
use BU_3VX2  BU_3VX2_30
timestamp 1529525674
transform -1 0 10584 0 -1 952
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_NO2_3VX4_1
timestamp 1529525674
transform 1 0 10584 0 -1 952
box 0 0 560 896
use NO2_3VX4  NO2_3VX4_1
timestamp 1529525674
transform 1 0 11144 0 -1 952
box 0 0 1344 896
use NA2I1_3VX2  NA2I1_3VX2_4
timestamp 1529525674
transform -1 0 13496 0 -1 952
box 0 0 1008 896
use NA2I1_3VX2  NA2I1_3VX2_1
timestamp 1529525674
transform 1 0 13496 0 -1 952
box 0 0 1008 896
use BU_3VX2  BU_3VX2_56
timestamp 1529525674
transform -1 0 15176 0 -1 952
box 0 0 672 896
use OR4_3VX1  OR4_3VX1_2
timestamp 1529525674
transform 1 0 15176 0 -1 952
box 0 0 1232 896
use IN_3VX0  IN_3VX0_3
timestamp 1529525674
transform -1 0 16744 0 -1 952
box 0 0 336 896
use DECAP7_3V  DECAP7_3V_0_1_0
timestamp 1529525674
transform 1 0 16744 0 -1 952
box 0 0 784 896
use BU_3VX2  BU_3VX2_53
timestamp 1529525674
transform 1 0 17528 0 -1 952
box 0 0 672 896
use BU_3VX2  BU_3VX2_37
timestamp 1529525674
transform 1 0 18200 0 -1 952
box 0 0 672 896
use BU_3VX2  BU_3VX2_38
timestamp 1529525674
transform 1 0 18872 0 -1 952
box 0 0 672 896
use DECAP5_3V  DECAP5_3V_0_DFRRQ_3VX4_2
timestamp 1529525674
transform -1 0 20104 0 -1 952
box 0 0 560 896
use DFRRQ_3VX4  DFRRQ_3VX4_2
timestamp 1529525674
transform -1 0 23688 0 -1 952
box 0 0 3584 896
<< labels >>
rlabel metaltpl s 5992 -336 6776 56 8 vdd3
port 0 nsew
rlabel metaltpl s 16408 -336 17192 56 8 gnd
port 1 nsew
rlabel metal3 s -252 18676 -196 18732 4 RST
port 2 nsew
rlabel metal3 s -252 18452 -196 18508 4 SCK
port 3 nsew
rlabel metal3 s -252 18228 -196 18284 4 SDI
port 4 nsew
rlabel metal3 s -252 18004 -196 18060 4 CSB
port 5 nsew
rlabel metal3 s 24052 3108 24108 3164 6 trap
port 6 nsew
rlabel metal3 s 24052 15092 24108 15148 6 pass_thru_sdo
port 7 nsew
rlabel metal2 s 13076 20916 13132 20972 6 mask_rev_in[0]
port 8 nsew
rlabel metal2 s 21364 20916 21420 20972 6 mask_rev_in[1]
port 9 nsew
rlabel metal2 s 22484 20916 22540 20972 6 mask_rev_in[2]
port 10 nsew
rlabel metal2 s 22708 20916 22764 20972 6 mask_rev_in[3]
port 11 nsew
rlabel metal3 s -252 17780 -196 17836 4 SDO
port 12 nsew
rlabel metal3 s -252 17556 -196 17612 4 sdo_enb
port 13 nsew
rlabel metal3 s 24052 12404 24108 12460 6 xtal_ena
port 14 nsew
rlabel metal3 s 24052 4004 24108 4060 6 reg_ena
port 15 nsew
rlabel metal3 s 24052 11396 24108 11452 6 pll_vco_ena
port 16 nsew
rlabel metal3 s 24052 11172 24108 11228 6 pll_cp_ena
port 17 nsew
rlabel metal3 s 24052 6692 24108 6748 6 pll_bias_ena
port 18 nsew
rlabel metal2 s 18340 -252 18396 -196 8 pll_trim[0]
port 19 nsew
rlabel metal2 s 18564 -252 18620 -196 8 pll_trim[1]
port 20 nsew
rlabel metal2 s 19124 -252 19180 -196 8 pll_trim[2]
port 21 nsew
rlabel metal2 s 22148 -252 22204 -196 8 pll_trim[3]
port 22 nsew
rlabel metal3 s 24052 4900 24108 4956 6 pll_bypass
port 23 nsew
rlabel metal3 s 24052 12180 24108 12236 6 pll_vco_in
port 24 nsew
rlabel metal2 s 18116 -252 18172 -196 8 tm_nvcp[0]
port 25 nsew
rlabel metal2 s 17892 -252 17948 -196 8 tm_nvcp[1]
port 26 nsew
rlabel metal2 s 17668 -252 17724 -196 8 tm_nvcp[2]
port 27 nsew
rlabel metal2 s 14756 -252 14812 -196 8 tm_nvcp[3]
port 28 nsew
rlabel metal3 s 24052 1316 24108 1372 6 irq
port 29 nsew
rlabel metal3 s 24052 3332 24108 3388 6 reset
port 30 nsew
rlabel metal2 s 10164 -252 10220 -196 8 pass_thru_reset
port 31 nsew
rlabel metal3 s 24052 14868 24108 14924 6 pass_thru_sck
port 32 nsew
rlabel metal3 s 24052 14644 24108 14700 6 pass_thru_csb
port 33 nsew
rlabel metal3 s 24052 14420 24108 14476 6 pass_thru_sdi
port 34 nsew
rlabel metal3 s 24052 17780 24108 17836 6 mfgr_id[0]
port 35 nsew
rlabel metal3 s 24052 17556 24108 17612 6 mfgr_id[1]
port 36 nsew
rlabel metal3 s 24052 17332 24108 17388 6 mfgr_id[2]
port 37 nsew
rlabel metal3 s 24052 17108 24108 17164 6 mfgr_id[3]
port 38 nsew
rlabel metal3 s 24052 16884 24108 16940 6 mfgr_id[4]
port 39 nsew
rlabel metal3 s 24052 16660 24108 16716 6 mfgr_id[5]
port 40 nsew
rlabel metal3 s 24052 16436 24108 16492 6 mfgr_id[6]
port 41 nsew
rlabel metal3 s 24052 16212 24108 16268 6 mfgr_id[7]
port 42 nsew
rlabel metal3 s 24052 15988 24108 16044 6 mfgr_id[8]
port 43 nsew
rlabel metal3 s 24052 15764 24108 15820 6 mfgr_id[9]
port 44 nsew
rlabel metal3 s 24052 15540 24108 15596 6 mfgr_id[10]
port 45 nsew
rlabel metal3 s 24052 15316 24108 15372 6 mfgr_id[11]
port 46 nsew
rlabel metal3 s 24052 12628 24108 12684 6 prod_id[0]
port 47 nsew
rlabel metal3 s 24052 12852 24108 12908 6 prod_id[1]
port 48 nsew
rlabel metal3 s 24052 13076 24108 13132 6 prod_id[2]
port 49 nsew
rlabel metal3 s 24052 13300 24108 13356 6 prod_id[3]
port 50 nsew
rlabel metal3 s 24052 13524 24108 13580 6 prod_id[4]
port 51 nsew
rlabel metal3 s 24052 13748 24108 13804 6 prod_id[5]
port 52 nsew
rlabel metal3 s 24052 13972 24108 14028 6 prod_id[6]
port 53 nsew
rlabel metal3 s 24052 14196 24108 14252 6 prod_id[7]
port 54 nsew
rlabel metal3 s 24052 18676 24108 18732 6 mask_rev[0]
port 55 nsew
rlabel metal3 s 24052 18452 24108 18508 6 mask_rev[1]
port 56 nsew
rlabel metal3 s 24052 18228 24108 18284 6 mask_rev[2]
port 57 nsew
rlabel metal3 s 24052 18004 24108 18060 6 mask_rev[3]
port 58 nsew
<< end >>
