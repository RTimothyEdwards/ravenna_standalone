magic
tech EFXH018D
timestamp 1533305873
<< mimcap >>
rect -4445 4825 -2445 4840
rect -4445 2555 -4430 4825
rect -2460 2555 -2445 4825
rect -4445 2540 -2445 2555
rect -2180 4825 -180 4840
rect -2180 2555 -2165 4825
rect -195 2555 -180 4825
rect -2180 2540 -180 2555
rect 85 4825 2085 4840
rect 85 2555 100 4825
rect 2070 2555 2085 4825
rect 85 2540 2085 2555
rect 2350 4825 4350 4840
rect 2350 2555 2365 4825
rect 4335 2555 4350 4825
rect 2350 2540 4350 2555
rect -4445 2365 -2445 2380
rect -4445 95 -4430 2365
rect -2460 95 -2445 2365
rect -4445 80 -2445 95
rect -2180 2365 -180 2380
rect -2180 95 -2165 2365
rect -195 95 -180 2365
rect -2180 80 -180 95
rect 85 2365 2085 2380
rect 85 95 100 2365
rect 2070 95 2085 2365
rect 85 80 2085 95
rect 2350 2365 4350 2380
rect 2350 95 2365 2365
rect 4335 95 4350 2365
rect 2350 80 4350 95
rect -4445 -95 -2445 -80
rect -4445 -2365 -4430 -95
rect -2460 -2365 -2445 -95
rect -4445 -2380 -2445 -2365
rect -2180 -95 -180 -80
rect -2180 -2365 -2165 -95
rect -195 -2365 -180 -95
rect -2180 -2380 -180 -2365
rect 85 -95 2085 -80
rect 85 -2365 100 -95
rect 2070 -2365 2085 -95
rect 85 -2380 2085 -2365
rect 2350 -95 4350 -80
rect 2350 -2365 2365 -95
rect 4335 -2365 4350 -95
rect 2350 -2380 4350 -2365
rect -4445 -2555 -2445 -2540
rect -4445 -4825 -4430 -2555
rect -2460 -4825 -2445 -2555
rect -4445 -4840 -2445 -4825
rect -2180 -2555 -180 -2540
rect -2180 -4825 -2165 -2555
rect -195 -4825 -180 -2555
rect -2180 -4840 -180 -4825
rect 85 -2555 2085 -2540
rect 85 -4825 100 -2555
rect 2070 -4825 2085 -2555
rect 85 -4840 2085 -4825
rect 2350 -2555 4350 -2540
rect 2350 -4825 2365 -2555
rect 4335 -4825 4350 -2555
rect 2350 -4840 4350 -4825
<< mimcapcontact >>
rect -4430 2555 -2460 4825
rect -2165 2555 -195 4825
rect 100 2555 2070 4825
rect 2365 2555 4335 4825
rect -4430 95 -2460 2365
rect -2165 95 -195 2365
rect 100 95 2070 2365
rect 2365 95 4335 2365
rect -4430 -2365 -2460 -95
rect -2165 -2365 -195 -95
rect 100 -2365 2070 -95
rect 2365 -2365 4335 -95
rect -4430 -4825 -2460 -2555
rect -2165 -4825 -195 -2555
rect 100 -4825 2070 -2555
rect 2365 -4825 4335 -2555
<< metal4 >>
rect -4495 4876 -2300 4890
rect -4495 4840 -2360 4876
rect -4495 2540 -4445 4840
rect -2445 2540 -2360 4840
rect -4495 2504 -2360 2540
rect -2310 2504 -2300 4876
rect -4495 2490 -2300 2504
rect -2230 4876 -35 4890
rect -2230 4840 -95 4876
rect -2230 2540 -2180 4840
rect -180 2540 -95 4840
rect -2230 2504 -95 2540
rect -45 2504 -35 4876
rect -2230 2490 -35 2504
rect 35 4876 2230 4890
rect 35 4840 2170 4876
rect 35 2540 85 4840
rect 2085 2540 2170 4840
rect 35 2504 2170 2540
rect 2220 2504 2230 4876
rect 35 2490 2230 2504
rect 2300 4876 4495 4890
rect 2300 4840 4435 4876
rect 2300 2540 2350 4840
rect 4350 2540 4435 4840
rect 2300 2504 4435 2540
rect 4485 2504 4495 4876
rect 2300 2490 4495 2504
rect -4495 2416 -2300 2430
rect -4495 2380 -2360 2416
rect -4495 80 -4445 2380
rect -2445 80 -2360 2380
rect -4495 44 -2360 80
rect -2310 44 -2300 2416
rect -4495 30 -2300 44
rect -2230 2416 -35 2430
rect -2230 2380 -95 2416
rect -2230 80 -2180 2380
rect -180 80 -95 2380
rect -2230 44 -95 80
rect -45 44 -35 2416
rect -2230 30 -35 44
rect 35 2416 2230 2430
rect 35 2380 2170 2416
rect 35 80 85 2380
rect 2085 80 2170 2380
rect 35 44 2170 80
rect 2220 44 2230 2416
rect 35 30 2230 44
rect 2300 2416 4495 2430
rect 2300 2380 4435 2416
rect 2300 80 2350 2380
rect 4350 80 4435 2380
rect 2300 44 4435 80
rect 4485 44 4495 2416
rect 2300 30 4495 44
rect -4495 -44 -2300 -30
rect -4495 -80 -2360 -44
rect -4495 -2380 -4445 -80
rect -2445 -2380 -2360 -80
rect -4495 -2416 -2360 -2380
rect -2310 -2416 -2300 -44
rect -4495 -2430 -2300 -2416
rect -2230 -44 -35 -30
rect -2230 -80 -95 -44
rect -2230 -2380 -2180 -80
rect -180 -2380 -95 -80
rect -2230 -2416 -95 -2380
rect -45 -2416 -35 -44
rect -2230 -2430 -35 -2416
rect 35 -44 2230 -30
rect 35 -80 2170 -44
rect 35 -2380 85 -80
rect 2085 -2380 2170 -80
rect 35 -2416 2170 -2380
rect 2220 -2416 2230 -44
rect 35 -2430 2230 -2416
rect 2300 -44 4495 -30
rect 2300 -80 4435 -44
rect 2300 -2380 2350 -80
rect 4350 -2380 4435 -80
rect 2300 -2416 4435 -2380
rect 4485 -2416 4495 -44
rect 2300 -2430 4495 -2416
rect -4495 -2504 -2300 -2490
rect -4495 -2540 -2360 -2504
rect -4495 -4840 -4445 -2540
rect -2445 -4840 -2360 -2540
rect -4495 -4876 -2360 -4840
rect -2310 -4876 -2300 -2504
rect -4495 -4890 -2300 -4876
rect -2230 -2504 -35 -2490
rect -2230 -2540 -95 -2504
rect -2230 -4840 -2180 -2540
rect -180 -4840 -95 -2540
rect -2230 -4876 -95 -4840
rect -45 -4876 -35 -2504
rect -2230 -4890 -35 -4876
rect 35 -2504 2230 -2490
rect 35 -2540 2170 -2504
rect 35 -4840 85 -2540
rect 2085 -4840 2170 -2540
rect 35 -4876 2170 -4840
rect 2220 -4876 2230 -2504
rect 35 -4890 2230 -4876
rect 2300 -2504 4495 -2490
rect 2300 -2540 4435 -2504
rect 2300 -4840 2350 -2540
rect 4350 -4840 4435 -2540
rect 2300 -4876 4435 -4840
rect 4485 -4876 4495 -2504
rect 2300 -4890 4495 -4876
<< viatp >>
rect -2360 2504 -2310 4876
rect -95 2504 -45 4876
rect 2170 2504 2220 4876
rect 4435 2504 4485 4876
rect -2360 44 -2310 2416
rect -95 44 -45 2416
rect 2170 44 2220 2416
rect 4435 44 4485 2416
rect -2360 -2416 -2310 -44
rect -95 -2416 -45 -44
rect 2170 -2416 2220 -44
rect 4435 -2416 4485 -44
rect -2360 -4876 -2310 -2504
rect -95 -4876 -45 -2504
rect 2170 -4876 2220 -2504
rect 4435 -4876 4485 -2504
<< metaltp >>
rect -3480 4825 -3410 4920
rect -2370 4876 -2300 4920
rect -3480 2365 -3410 2555
rect -2370 2504 -2360 4876
rect -2310 2504 -2300 4876
rect -1215 4825 -1145 4920
rect -105 4876 -35 4920
rect -2370 2416 -2300 2504
rect -3480 -95 -3410 95
rect -2370 44 -2360 2416
rect -2310 44 -2300 2416
rect -1215 2365 -1145 2555
rect -105 2504 -95 4876
rect -45 2504 -35 4876
rect 1050 4825 1120 4920
rect 2160 4876 2230 4920
rect -105 2416 -35 2504
rect -2370 -44 -2300 44
rect -3480 -2555 -3410 -2365
rect -2370 -2416 -2360 -44
rect -2310 -2416 -2300 -44
rect -1215 -95 -1145 95
rect -105 44 -95 2416
rect -45 44 -35 2416
rect 1050 2365 1120 2555
rect 2160 2504 2170 4876
rect 2220 2504 2230 4876
rect 3315 4825 3385 4920
rect 4425 4876 4495 4920
rect 2160 2416 2230 2504
rect -105 -44 -35 44
rect -2370 -2504 -2300 -2416
rect -3480 -4920 -3410 -4825
rect -2370 -4876 -2360 -2504
rect -2310 -4876 -2300 -2504
rect -1215 -2555 -1145 -2365
rect -105 -2416 -95 -44
rect -45 -2416 -35 -44
rect 1050 -95 1120 95
rect 2160 44 2170 2416
rect 2220 44 2230 2416
rect 3315 2365 3385 2555
rect 4425 2504 4435 4876
rect 4485 2504 4495 4876
rect 4425 2416 4495 2504
rect 2160 -44 2230 44
rect -105 -2504 -35 -2416
rect -2370 -4920 -2300 -4876
rect -1215 -4920 -1145 -4825
rect -105 -4876 -95 -2504
rect -45 -4876 -35 -2504
rect 1050 -2555 1120 -2365
rect 2160 -2416 2170 -44
rect 2220 -2416 2230 -44
rect 3315 -95 3385 95
rect 4425 44 4435 2416
rect 4485 44 4495 2416
rect 4425 -44 4495 44
rect 2160 -2504 2230 -2416
rect -105 -4920 -35 -4876
rect 1050 -4920 1120 -4825
rect 2160 -4876 2170 -2504
rect 2220 -4876 2230 -2504
rect 3315 -2555 3385 -2365
rect 4425 -2416 4435 -44
rect 4485 -2416 4495 -44
rect 4425 -2504 4495 -2416
rect 2160 -4920 2230 -4876
rect 3315 -4920 3385 -4825
rect 4425 -4876 4435 -2504
rect 4485 -4876 4495 -2504
rect 4425 -4920 4495 -4876
<< boundary >>
rect -4495 2490 -2395 4890
rect -2230 2490 -130 4890
rect 35 2490 2135 4890
rect 2300 2490 4400 4890
rect -4495 30 -2395 2430
rect -2230 30 -130 2430
rect 35 30 2135 2430
rect 2300 30 4400 2430
rect -4495 -2430 -2395 -30
rect -2230 -2430 -130 -30
rect 35 -2430 2135 -30
rect 2300 -2430 4400 -30
rect -4495 -4890 -2395 -2490
rect -2230 -4890 -130 -2490
rect 35 -4890 2135 -2490
rect 2300 -4890 4400 -2490
<< properties >>
string parameters w 20.00 l 23.00 val 474.62 carea 1.00 cperi 0.17 nx 4 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
