magic
tech EFXH018D
magscale 1 2
timestamp 1523029302
<< metal2 >>
tri 9 1739 217 1947 se
rect 217 1739 857 1947
tri 857 1739 1065 1947 sw
rect 9 1723 1065 1739
rect 9 1105 217 1723
tri 217 1611 329 1723 nw
tri 745 1611 857 1723 ne
tri 217 1105 329 1217 sw
tri 745 1105 857 1217 se
rect 857 1105 1065 1723
tri 9 1001 113 1105 ne
tri 9 897 113 1001 se
rect 113 897 961 1105
tri 961 1001 1065 1105 nw
tri 961 897 1065 1001 sw
rect 9 235 217 897
tri 217 785 329 897 nw
tri 745 785 857 897 ne
tri 217 235 329 347 sw
tri 745 235 857 347 se
rect 857 235 1065 897
tri 9 27 217 235 ne
rect 217 27 857 235
tri 857 27 1065 235 nw
<< end >>
