magic
tech EFXH018D
magscale 1 2
timestamp 1555546887
<< error_s >>
rect -89573 313552 -89173 320352
rect -85573 313552 -85173 320352
rect -68773 313552 -68373 320352
rect -51973 313552 -51573 320352
rect -35273 313552 -34773 320352
rect 112627 313552 113127 320352
rect 129427 313552 129827 320352
rect 146227 313552 146627 320352
rect 163027 313552 163427 320352
rect 179827 313552 180227 320352
rect 196627 313552 197027 320352
rect 213427 313552 213827 320352
rect 230227 313552 230627 320352
rect 234227 313552 234627 320352
rect 30829 309039 32000 309067
rect -28933 308171 -25353 308199
rect -28933 303753 -28905 308171
rect -25381 303753 -25353 308171
rect 9947 307753 13287 307781
rect 9947 303932 9975 307753
rect 13259 303932 13287 307753
rect 9947 303904 13287 303932
rect -28933 303725 -25353 303753
rect 30829 302696 30857 309039
rect 97101 308771 101491 308799
rect 97101 302696 97129 308771
rect 101463 302696 101491 308771
rect 30829 302668 32000 302696
rect 97101 302668 101491 302696
rect -89573 291928 -89173 298328
rect -85573 291928 -85173 298328
rect -68773 291928 -68373 298328
rect -51973 291928 -51573 298328
rect -35273 291928 -34773 298328
rect 112627 291928 113127 298328
rect 129427 291928 129827 298328
rect 146227 291928 146627 298328
rect 163027 291928 163427 298328
rect 179827 291928 180227 298328
rect 196627 291928 197027 298328
rect 213427 291928 213827 298328
rect 230227 291928 230627 298328
rect 234227 291928 234627 298328
rect -89773 290700 -89173 291428
rect -85773 290700 -85173 291428
rect -68973 290700 -68373 291428
rect -52173 290700 -51573 291428
rect -35373 290700 -34773 291428
rect 112527 290700 113127 291428
rect 129227 290700 129827 291428
rect 146027 290700 146627 291428
rect 162827 290700 163427 291428
rect 179627 290700 180227 291428
rect 196427 290700 197027 291428
rect 213227 290700 213827 291428
rect 230027 290700 230627 291428
rect 234027 290700 234627 291428
rect -89773 289600 -89173 290200
rect -85773 289600 -85173 290200
rect -68973 289600 -68373 290200
rect -52173 289600 -51573 290200
rect -35373 289600 -34773 290200
rect 112527 289600 113127 290200
rect 129227 289600 129827 290200
rect 146027 289600 146627 290200
rect 162827 289600 163427 290200
rect 179627 289600 180227 290200
rect 196427 289600 197027 290200
rect 213227 289600 213827 290200
rect 230027 289600 230627 290200
rect 234027 289600 234627 290200
rect -89773 288500 -89173 289100
rect -85773 288500 -85173 289100
rect -68973 288500 -68373 289100
rect -52173 288500 -51573 289100
rect -35373 288500 -34773 289100
rect 112527 288500 113127 289100
rect 129227 288500 129827 289100
rect 146027 288500 146627 289100
rect 162827 288500 163427 289100
rect 179627 288500 180227 289100
rect 196427 288500 197027 289100
rect 213227 288500 213827 289100
rect 230027 288500 230627 289100
rect 234027 288852 234627 289100
rect 234027 288500 234875 288852
rect -91521 287852 -90921 288452
rect -90421 287852 -89821 288452
rect 234275 288252 234875 288500
rect 235375 288252 235975 288852
rect 236475 288252 237203 288852
rect 237703 288452 244103 288852
rect 259327 288452 266127 288852
rect 234275 284352 234875 284952
rect 235375 284352 235975 284952
rect 236475 284352 237203 284952
rect 237703 284452 244103 284952
rect 259327 284452 266127 284952
rect 248443 273288 254574 273316
rect -121673 271252 -114873 271652
rect -99649 271252 -93249 271652
rect -92749 271052 -92021 271652
rect -91521 271052 -90921 271652
rect -90421 271052 -89821 271652
rect 195387 268952 195447 269012
rect 248443 268954 248471 273288
rect 254546 268954 254574 273288
rect 248443 268926 254574 268954
rect 195387 268792 195447 268852
rect -91521 253852 -90921 254452
rect -90421 253852 -89821 254452
rect -121673 252052 -114873 252452
rect -99649 252052 -93249 252452
rect -92749 251852 -92021 252452
rect -91521 251852 -90921 252452
rect -90421 251852 -89821 252452
rect -121673 248052 -114873 248452
rect -99649 248052 -93249 248452
rect -92749 247852 -92021 248452
rect -91521 247852 -90921 248452
rect -90421 247852 -89821 248452
rect -121673 231252 -114873 231652
rect -99649 231252 -93249 231652
rect -92749 231052 -92021 231652
rect -91521 231052 -90921 231652
rect -90421 231052 -89821 231652
rect -121673 214452 -114873 214852
rect -99649 214452 -93249 214852
rect -92749 214252 -92021 214852
rect -91521 214252 -90921 214852
rect -90421 214252 -89821 214852
rect 248443 207150 254842 207178
rect 248443 202682 248471 207150
rect 254814 202682 254842 207150
rect 248443 202654 254842 202682
rect -121673 197652 -114873 198052
rect -99649 197652 -93249 198052
rect -92749 197452 -92021 198052
rect -91521 197452 -90921 198052
rect -90421 197452 -89821 198052
rect 234275 191652 234875 192252
rect 235375 191652 235975 192252
rect 236475 191652 237203 192252
rect 237703 191752 244103 192252
rect 259327 191752 266127 192252
rect 234275 181652 234875 182252
rect 235375 181652 235975 182252
rect 236475 181652 237203 182252
rect 237703 181852 244103 182252
rect 259327 181852 266127 182252
rect -121673 180852 -114873 181252
rect -99649 180852 -93249 181252
rect -92749 180652 -92021 181252
rect -91521 180652 -90921 181252
rect -90421 180652 -89821 181252
rect 234275 164852 234875 165452
rect 235375 164852 235975 165452
rect 236475 164852 237203 165452
rect 237703 165052 244103 165452
rect 259327 165052 266127 165452
rect -121673 164052 -114873 164452
rect -99649 164052 -93249 164452
rect -92749 163852 -92021 164452
rect -91521 163852 -90921 164452
rect -90421 163852 -89821 164452
rect 234275 160852 234875 161452
rect 235375 160852 235975 161452
rect 236475 160852 237203 161452
rect 237703 161052 244103 161452
rect 259327 161052 266127 161452
rect -121673 147252 -114873 147652
rect -99649 147252 -93249 147652
rect -92749 147052 -92021 147652
rect -91521 147052 -90921 147652
rect -90421 147052 -89821 147652
rect 234275 144052 234875 144652
rect 235375 144052 235975 144652
rect 236475 144052 237203 144652
rect 237703 144252 244103 144652
rect 259327 144252 266127 144652
rect -121673 130452 -114873 130852
rect -99649 130452 -93249 130852
rect -92749 130252 -92021 130852
rect -91521 130252 -90921 130852
rect -90421 130252 -89821 130852
rect 234275 127252 234875 127852
rect 235375 127252 235975 127852
rect 236475 127252 237203 127852
rect 237703 127452 244103 127852
rect 259327 127452 266127 127852
rect -121673 113652 -114873 114052
rect -99649 113652 -93249 114052
rect -92749 113452 -92021 114052
rect -91521 113452 -90921 114052
rect -90421 113452 -89821 114052
rect 234275 110452 234875 111052
rect 235375 110452 235975 111052
rect 236475 110452 237203 111052
rect 237703 110652 244103 111052
rect 259327 110652 266127 111052
rect 234275 100452 234875 101052
rect 235375 100452 235975 101052
rect 236475 100452 237203 101052
rect 237703 100652 244103 101052
rect 259327 100652 266127 101052
rect -121673 96852 -114873 97252
rect -99649 96852 -93249 97252
rect -92749 96652 -92021 97252
rect -91521 96652 -90921 97252
rect -90421 96652 -89821 97252
rect 234275 83652 234875 84252
rect 235375 83652 235975 84252
rect 236475 83652 237203 84252
rect 237703 83852 244103 84252
rect 259327 83852 266127 84252
rect -121673 80052 -114873 80452
rect -99649 80052 -93249 80452
rect -92749 79852 -92021 80452
rect -91521 79852 -90921 80452
rect -90421 79852 -89821 80452
rect 284228 68282 284828 68882
rect 285328 68282 285928 68882
rect 286428 68382 287156 68882
rect 287656 68382 288000 68882
rect 286428 68282 287311 68382
rect 234275 66852 234875 67452
rect 235375 66852 235975 67452
rect 236475 66852 237203 67452
rect 237703 67052 244103 67452
rect 259327 67052 266127 67452
rect -121673 63252 -114873 63652
rect -99649 63252 -93249 63652
rect -92749 63052 -92021 63652
rect -91521 63052 -90921 63652
rect -90421 63052 -89821 63652
rect -171892 61892 -165092 62292
rect -149868 61892 -143468 62292
rect -142968 61692 -142240 62292
rect -141740 61692 -141140 62292
rect -140640 61692 -140040 62292
rect 284228 51482 284828 52082
rect 285328 51482 285928 52082
rect 286428 51482 287156 52082
rect 287656 51682 294056 52082
rect 309280 51682 316080 52082
rect 234275 50052 234875 50652
rect 235375 50052 235975 50652
rect 236475 50052 237203 50652
rect 237703 50252 244103 50652
rect 259327 50252 266127 50652
rect -121673 46452 -114873 46652
rect -99649 46452 -93249 46652
rect -92749 46052 -92021 46652
rect -91521 46052 -90921 46652
rect -90421 46052 -89821 46652
rect -171892 45092 -165092 45592
rect -149868 45092 -143468 45592
rect -142968 45092 -142240 45592
rect -143123 44992 -142240 45092
rect -141740 44992 -141140 45592
rect -140640 44992 -140040 45592
rect 284228 34682 284828 35282
rect 285328 34682 285928 35282
rect 286428 34682 287156 35282
rect 287656 34882 294056 35282
rect 309280 34882 316080 35282
rect 234275 33252 234875 33852
rect 235375 33252 235975 33852
rect 236475 33252 237203 33852
rect 237703 33452 244103 33852
rect 259327 33452 266127 33852
rect -121673 29452 -114873 29852
rect -99649 29452 -93249 29852
rect -92749 29252 -92021 29852
rect -91521 29252 -90921 29852
rect -90421 29252 -89821 29852
rect 284228 17882 284828 18482
rect 285328 17882 285928 18482
rect 286428 17882 287156 18482
rect 287656 18082 294056 18482
rect 309280 18082 316080 18482
rect 234275 16452 234875 17052
rect 235375 16452 235975 17052
rect 236475 16452 237203 17052
rect 237703 16652 244103 17052
rect 259327 16652 266127 17052
rect -121673 12652 -114873 13052
rect -99649 12652 -93249 13052
rect -92749 12452 -92021 13052
rect -91521 12452 -90921 13052
rect -90421 12452 -89821 13052
rect 234275 12452 234875 13052
rect 235375 12452 235975 13052
rect 236475 12452 237203 13052
rect 237703 12652 244103 13052
rect 259327 12652 266127 13052
rect -89773 11804 -89173 12404
rect -85773 11804 -85173 12404
rect -68973 11804 -68373 12404
rect -52173 11804 -51573 12404
rect -48173 11804 -47573 12404
rect -47073 11804 -46473 12404
rect -30373 11804 -29773 12404
rect -26373 11804 -25773 12404
rect -9573 11804 -8973 12404
rect 7227 11804 7827 12404
rect 24027 11804 24627 12404
rect 40827 11804 41427 12404
rect 41927 11804 42527 12404
rect 49827 11804 50427 12404
rect 66627 11804 67227 12404
rect 83427 11804 84027 12404
rect 100227 11804 100827 12404
rect 117027 11804 117627 12404
rect 133827 11804 134427 12404
rect 150627 11804 151227 12404
rect 167427 11804 168027 12404
rect 184227 11804 184827 12404
rect 201027 11804 201627 12404
rect 217827 11804 218427 12404
rect 227827 11804 228427 12404
rect 231827 11804 232427 12404
rect 233827 11804 234427 12404
rect -89773 10704 -89173 11304
rect -85773 10704 -85173 11304
rect -68973 10704 -68373 11304
rect -52173 10704 -51573 11304
rect -48173 10704 -47573 11304
rect -47073 10704 -46473 11304
rect -30373 10704 -29773 11304
rect -26373 10704 -25773 11304
rect -9573 10704 -8973 11304
rect 7227 10704 7827 11304
rect 24027 10704 24627 11304
rect 40827 10704 41427 11304
rect 41927 10704 42527 11304
rect 49827 10704 50427 11304
rect 66627 10704 67227 11304
rect 83427 10704 84027 11304
rect 100227 10704 100827 11304
rect 117027 10704 117627 11304
rect 133827 10704 134427 11304
rect 150627 10704 151227 11304
rect 167427 10704 168027 11304
rect 184227 10704 184827 11304
rect 201027 10704 201627 11304
rect 217827 10704 218427 11304
rect 227827 10704 228427 11304
rect 231827 10704 232427 11304
rect 233827 10704 234427 11304
rect -89773 9476 -89173 10204
rect -85773 9476 -85173 10204
rect -68973 9476 -68373 10204
rect -52173 9476 -51573 10204
rect -48173 9476 -47573 10204
rect -47073 9476 -46473 10204
rect -30373 9476 -29773 10204
rect -26373 9476 -25773 10204
rect -9573 9476 -8973 10204
rect 7227 9476 7827 10204
rect 24027 9476 24627 10204
rect 40827 9476 41427 10204
rect 41927 9476 42527 10204
rect 49827 9476 50427 10204
rect 66627 9476 67227 10204
rect 83427 9476 84027 10204
rect 100227 9476 100827 10204
rect 117027 9476 117627 10204
rect 133827 9476 134427 10204
rect 150627 9476 151227 10204
rect 167427 9476 168027 10204
rect 184227 9476 184827 10204
rect 201027 9476 201627 10204
rect 217827 9476 218427 10204
rect 227827 9476 228427 10204
rect 231827 9476 232427 10204
rect 233827 9476 234427 10204
rect -89573 2576 -89173 8976
rect -85573 2576 -85173 8976
rect -68773 2576 -68373 8976
rect -51973 2576 -51573 8976
rect -48073 2576 -47573 8976
rect -46973 2576 -46473 8976
rect -30173 2576 -29773 8976
rect -26173 2576 -25773 8976
rect -9373 2576 -8973 8976
rect 7427 2576 7827 8976
rect 24227 2576 24627 8976
rect 40927 2576 41427 8976
rect 42027 2576 42527 8976
rect 50027 2576 50427 8976
rect 66827 2576 67227 8976
rect 83627 2576 84027 8976
rect 100427 2576 100827 8976
rect 117227 2576 117627 8976
rect 134027 2576 134427 8976
rect 150827 2576 151227 8976
rect 167627 2576 168027 8976
rect 184427 2576 184827 8976
rect 201227 2576 201627 8976
rect 218027 2576 218427 8976
rect 228027 2576 228427 8976
rect 232027 2576 232427 8976
rect 234227 2576 234427 8976
rect 284228 1182 284828 1782
rect 285328 1182 285928 1782
rect 286428 1282 287156 1782
rect 287656 1282 294056 1782
rect 309280 1282 316080 1782
rect 286428 1182 287311 1282
rect -89573 -19448 -89173 -12648
rect -85573 -19448 -85173 -12648
rect -68773 -19448 -68373 -12648
rect -51973 -19448 -51573 -12648
rect -48073 -19448 -47573 -12648
rect -46973 -19448 -46473 -12648
rect -30173 -19448 -29773 -12648
rect -26173 -19448 -25773 -12648
rect -9373 -19448 -8973 -12648
rect 7427 -19448 7827 -12648
rect 24227 -19448 24627 -12648
rect 40927 -19448 41427 -12648
rect 42027 -19448 42527 -12648
rect 50027 -19448 50427 -12648
rect 66827 -19448 67227 -12648
rect 83627 -19448 84027 -12648
rect 100427 -19448 100827 -12648
rect 117227 -19448 117627 -12648
rect 134027 -19448 134427 -12648
rect 150827 -19448 151227 -12648
rect 167627 -19448 168027 -12648
rect 184427 -19448 184827 -12648
rect 201227 -19448 201627 -12648
rect 218027 -19448 218427 -12648
rect 228027 -19448 228427 -12648
rect 232027 -19448 232427 -12648
rect 234227 -19448 234427 -12648
<< metal1 >>
rect -80670 301781 -73670 308781
rect -63870 301781 -56870 308781
rect -47070 301781 -40070 308781
rect 151388 302860 158388 309860
rect 168188 302860 175188 309860
rect 184445 303090 191445 310090
rect 201619 303242 208619 310242
rect 218945 302940 225945 309940
rect -110746 236073 -103746 243073
rect -110746 219273 -103746 226273
rect -110746 202473 -103746 209473
rect -110746 185673 -103746 192673
rect -110746 168873 -103746 175873
rect -110746 152073 -103746 159073
rect 247838 149085 254838 156085
rect -110746 135273 -103746 142273
rect 247838 132285 254838 139285
rect -110746 118473 -103746 125473
rect 247838 115485 254838 122485
rect -110746 101673 -103746 108673
rect -110746 84873 -103746 91873
rect 247838 88685 254838 95685
rect -110746 68073 -103746 75073
rect 247838 71885 254838 78885
rect -110746 51273 -103746 58273
rect 247838 55085 254838 62085
rect 247838 38285 254838 45285
rect 247838 21485 254838 28485
rect -64077 -8451 -57077 -1451
rect -42277 -8451 -35277 -1451
rect -21477 -8451 -14477 -1451
rect -4677 -8451 2323 -1451
rect 12123 -8451 19123 -1451
rect 54723 -8451 61723 -1451
rect 71523 -8451 78523 -1451
rect 88323 -8451 95323 -1451
rect 105123 -8451 112123 -1451
rect 121923 -8451 128923 -1451
rect 138723 -8451 145723 -1451
rect 155523 -8451 162523 -1451
<< metaltpl >>
rect -28441 304587 -25963 307436
rect 10336 304449 12814 307298
use CORNERESDF  CORNERESDF_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -121673 -1 0 320352
box 0 0 32000 32000
use FILLER20F  FILLER20F_3 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform -1 0 -85673 0 -1 320352
box 0 0 4000 32000
use BBCUD4F  BBCUD4F_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform -1 0 -68873 0 -1 320352
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_0
timestamp 1529526440
transform -1 0 -52073 0 -1 320352
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_1
timestamp 1529526440
transform -1 0 -35273 0 -1 320352
box 0 0 16800 32000
use axtoc02_3v3  axtoc02_3v3_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1516677002
transform -1 0 19927 0 -1 320352
box 0 0 55200 31882
use FILLER02F  FILLER02F_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -121673 -1 0 288352
box 0 0 400 32000
use GNDORPADF  GNDORPADF_7 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -121673 -1 0 287952
box 0 0 16800 32000
use VDDORPADF  VDDORPADF_3 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -121673 -1 0 271152
box 0 0 16800 32000
use FILLER02F  FILLER02F_0
timestamp 1529526440
transform 0 1 -121673 -1 0 254352
box 0 0 400 32000
use FILLER10F  FILLER10F_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -121673 -1 0 253952
box 0 0 2000 32000
use FILLER20F  FILLER20F_5
timestamp 1529526440
transform 0 1 -121673 -1 0 251952
box 0 0 4000 32000
use aregc01_3v3  aregc01_3v3_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1516677094
transform -1 0 112527 0 -1 320352
box 0 0 92600 70740
use GNDORPADF  GNDORPADF_1
timestamp 1529526440
transform -1 0 129327 0 -1 320352
box 0 0 16800 32000
use VDDORPADF  VDDORPADF_1
timestamp 1529526440
transform -1 0 146127 0 -1 320352
box 0 0 16800 32000
use APR00DF  APR00DF_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform -1 0 162927 0 -1 320352
box 0 0 16800 32000
use APR00DF  APR00DF_1
timestamp 1529526440
transform -1 0 179727 0 -1 320352
box 0 0 16800 32000
use APR00DF  APR00DF_2
timestamp 1529526440
transform -1 0 196527 0 -1 320352
box 0 0 16800 32000
use APR00DF  APR00DF_3
timestamp 1529526440
transform -1 0 213327 0 -1 320352
box 0 0 16800 32000
use APR00DF  APR00DF_4
timestamp 1529526440
transform -1 0 230127 0 -1 320352
box 0 0 16800 32000
use FILLER20F  FILLER20F_2
timestamp 1529526440
transform 1 0 230127 0 -1 320352
box 0 0 4000 32000
use CORNERESDF  CORNERESDF_0
timestamp 1529526440
transform -1 0 266127 0 -1 320352
box 0 0 32000 32000
use FILLER20F  FILLER20F_4
timestamp 1529526440
transform 0 -1 266127 -1 0 288352
box 0 0 4000 32000
use BBCUD4F  BBCUD4F_3
timestamp 1529526440
transform 0 1 -121673 -1 0 247952
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_4
timestamp 1529526440
transform 0 1 -121673 -1 0 231152
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_5
timestamp 1529526440
transform 0 1 -121673 -1 0 214352
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_6
timestamp 1529526440
transform 0 1 -121673 -1 0 197552
box 0 0 16800 32000
use aregc01_3v3  aregc01_3v3_1
timestamp 1516677094
transform 0 -1 266127 -1 0 284352
box 0 0 92600 70740
use BBCUD4F  BBCUD4F_7
timestamp 1529526440
transform 0 1 -121673 -1 0 180752
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_8
timestamp 1529526440
transform 0 1 -121673 -1 0 163952
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_9
timestamp 1529526440
transform 0 1 -121673 -1 0 147152
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_10
timestamp 1529526440
transform 0 1 -121673 -1 0 130352
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_11
timestamp 1529526440
transform 0 1 -121673 -1 0 113552
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_12
timestamp 1529526440
transform 0 1 -121673 -1 0 96752
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_16
timestamp 1529526440
transform 0 1 -171892 -1 0 78592
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_17
timestamp 1529526440
transform 0 1 -171892 -1 0 61792
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_13
timestamp 1529526440
transform 0 1 -121673 -1 0 79952
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_14
timestamp 1529526440
transform 0 1 -121673 -1 0 63152
box 0 0 16800 32000
use FILLER01F  FILLER01F_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -121673 -1 0 46352
box 0 0 200 32000
use VDDORPADF  VDDORPADF_2
timestamp 1529526440
transform 0 1 -121673 -1 0 46152
box 0 0 16800 32000
use GNDORPADF  GNDORPADF_6
timestamp 1529526440
transform 0 1 -121673 -1 0 29352
box 0 0 16800 32000
use FILLER50F  FILLER50F_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 -1 266127 -1 0 191752
box 0 0 10000 32000
use GNDORPADF  GNDORPADF_2
timestamp 1529526440
transform 0 -1 266127 1 0 164952
box 0 0 16800 32000
use FILLER20F  FILLER20F_6
timestamp 1529526440
transform 0 -1 266127 1 0 160952
box 0 0 4000 32000
use VDDPADF  VDDPADF_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 -1 266127 1 0 144152
box 0 0 16800 32000
use VDDORPADF  VDDORPADF_0
timestamp 1529526440
transform 0 -1 266127 1 0 127352
box 0 0 16800 32000
use GNDORPADF  GNDORPADF_0
timestamp 1529526440
transform 0 -1 266127 1 0 110552
box 0 0 16800 32000
use FILLER50F  FILLER50F_1
timestamp 1529526440
transform 0 -1 266127 1 0 100552
box 0 0 10000 32000
use APR00DF  APR00DF_5
timestamp 1529526440
transform 0 -1 266127 1 0 83752
box 0 0 16800 32000
use APR00DF  APR00DF_6
timestamp 1529526440
transform 0 -1 266127 1 0 66952
box 0 0 16800 32000
use ICF  ICF_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 -1 266127 1 0 50152
box 0 0 16800 32000
use BT4F  BT4F_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 -1 266127 1 0 33352
box 0 0 16800 32000
use ICF  ICF_0
timestamp 1529526440
transform 0 -1 266127 1 0 16552
box 0 0 16800 32000
use FILLER20F  FILLER20F_7
timestamp 1529526440
transform 0 -1 266127 1 0 12552
box 0 0 4000 32000
use CORNERESDF  CORNERESDF_2
timestamp 1529526440
transform 1 0 -121673 0 1 -19448
box 0 0 32000 32000
use FILLER20F  FILLER20F_0
timestamp 1529526440
transform 1 0 -89673 0 1 -19448
box 0 0 4000 32000
use GNDORPADF  GNDORPADF_5
timestamp 1529526440
transform 1 0 -85673 0 1 -19448
box 0 0 16800 32000
use BBCUD4F  BBCUD4F_15
timestamp 1529526440
transform 1 0 -68873 0 1 -19448
box 0 0 16800 32000
use FILLER20F  FILLER20F_8
timestamp 1529526440
transform 1 0 -52073 0 1 -19448
box 0 0 4000 32000
use POWERCUTVDD3FC  POWERCUTVDD3FC_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_FC3V
timestamp 1516645956
transform -1 0 -47073 0 1 -19448
box 0 0 1000 32000
use ICFC  ICFC_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_FC3V
timestamp 1529532354
transform 1 0 -47073 0 1 -19448
box 0 0 16800 32000
use FILLER20FC  FILLER20FC_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_FC3V
timestamp 1529532354
transform 1 0 -30273 0 1 -19448
box 0 0 4000 32000
use ICFC  ICFC_1
timestamp 1529532354
transform 1 0 -26273 0 1 -19448
box 0 0 16800 32000
use ICFC  ICFC_2
timestamp 1529532354
transform 1 0 -9473 0 1 -19448
box 0 0 16800 32000
use BT4FC  BT4FC_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_FC3V
timestamp 1529532354
transform 1 0 7327 0 1 -19448
box 0 0 16800 32000
use VDDPADFC  VDDPADFC_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_FC3V
timestamp 1529532354
transform 1 0 24127 0 1 -19448
box 0 0 16800 32000
use POWERCUTVDD3FC  POWERCUTVDD3FC_1
timestamp 1516645956
transform 1 0 40927 0 1 -19448
box 0 0 1000 32000
use FILLER40F  FILLER40F_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 1 0 41927 0 1 -19448
box 0 0 8000 32000
use BBC4F  BBC4F_2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 1 0 49927 0 1 -19448
box 0 0 16800 32000
use BBC4F  BBC4F_3
timestamp 1529526440
transform 1 0 66727 0 1 -19448
box 0 0 16800 32000
use BBC4F  BBC4F_1
timestamp 1529526440
transform 1 0 83527 0 1 -19448
box 0 0 16800 32000
use BBC4F  BBC4F_0
timestamp 1529526440
transform 1 0 100327 0 1 -19448
box 0 0 16800 32000
use BT4F  BT4F_2
timestamp 1529526440
transform 1 0 117127 0 1 -19448
box 0 0 16800 32000
use BT4F  BT4F_1
timestamp 1529526440
transform 1 0 133927 0 1 -19448
box 0 0 16800 32000
use ICF  ICF_2
timestamp 1529526440
transform 1 0 150727 0 1 -19448
box 0 0 16800 32000
use GNDORPADF  GNDORPADF_3
timestamp 1529526440
transform 1 0 167527 0 1 -19448
box 0 0 16800 32000
use VDDORPADF  VDDORPADF_4
timestamp 1529526440
transform 1 0 184327 0 1 -19448
box 0 0 16800 32000
use VDDPADF  VDDPADF_1
timestamp 1529526440
transform 1 0 201127 0 1 -19448
box 0 0 16800 32000
use FILLER50F  FILLER50F_2
timestamp 1529526440
transform 1 0 217927 0 1 -19448
box 0 0 10000 32000
use FILLER20F  FILLER20F_1
timestamp 1529526440
transform 1 0 227927 0 1 -19448
box 0 0 4000 32000
use FILLER10F  FILLER10F_1
timestamp 1529526440
transform 1 0 231927 0 1 -19448
box 0 0 2000 32000
use FILLER01F  FILLER01F_1
timestamp 1529526440
transform 1 0 233927 0 1 -19448
box 0 0 200 32000
use CORNERESDF  CORNERESDF_3
timestamp 1529526440
transform 0 -1 266127 1 0 -19448
box 0 0 32000 32000
use ICF  ICF_3
timestamp 1529526440
transform 0 -1 316080 1 0 51582
box 0 0 16800 32000
use BT4F  BT4F_3
timestamp 1529526440
transform 0 -1 316080 1 0 34782
box 0 0 16800 32000
use BT4F  BT4F_4
timestamp 1529526440
transform 0 -1 316080 1 0 17982
box 0 0 16800 32000
use BT4F  BT4F_5
timestamp 1529526440
transform 0 -1 316080 1 0 1182
box 0 0 16800 32000
<< labels >>
rlabel metal1 -64077 -8451 -57077 -1451 0 gpio<15>
rlabel metal1 121923 -8451 128923 -1451 0 flash_csb
rlabel metal1 138723 -8451 145723 -1451 0 flash_clk
rlabel metal1 155523 -8451 162523 -1451 0 XCLK
rlabel metal1 -42277 -8451 -35277 -1451 0 SDI
rlabel metal1 12123 -8451 19123 -1451 0 SDO
rlabel metal1 -4677 -8451 2323 -1451 0 SCK
rlabel metal1 -21477 -8451 -14477 -1451 0 CSB
rlabel metal1 105123 -8451 112123 -1451 0 flash_io0
rlabel metal1 54723 -8451 61723 -1451 0 flash_io3
rlabel metal1 88323 -8451 95323 -1451 0 flash_io1
rlabel metal1 71523 -8451 78523 -1451 0 flash_io2
rlabel metal1 -47070 301781 -40070 308781 0 gpio<0>
rlabel metal1 -63870 301781 -56870 308781 0 gpio<1>
rlabel metal1 -80670 301781 -73670 308781 0 gpio<2>
rlabel metaltpl -28441 304587 -25963 307436 0 XO
rlabel metaltpl 10336 304449 12814 307298 0 XI
rlabel metal1 247838 21485 254838 28485 0 ser_rx
rlabel metal1 247838 38285 254838 45285 0 ser_tx
rlabel metal1 247838 115485 254838 122485 0 VSS
rlabel metal1 247838 55085 254838 62085 0 irq
rlabel metal1 247838 132285 254838 139285 0 VDD3V3
rlabel metal1 247838 149085 254838 156085 0 VDD1V8
rlabel metal1 -110746 236073 -103746 243073 0 gpio<3>
rlabel metal1 -110746 219273 -103746 226273 0 gpio<4>
rlabel metal1 -110746 202473 -103746 209473 0 gpio<5>
rlabel metal1 -110746 185673 -103746 192673 0 gpio<6>
rlabel metal1 -110746 168873 -103746 175873 0 gpio<7>
rlabel metal1 -110746 152073 -103746 159073 0 gpio<8>
rlabel metal1 -110746 135273 -103746 142273 0 gpio<9>
rlabel metal1 -110746 118473 -103746 125473 0 gpio<10>
rlabel metal1 -110746 101673 -103746 108673 0 gpio<11>
rlabel metal1 -110746 84873 -103746 91873 0 gpio<12>
rlabel metal1 -110746 68073 -103746 75073 0 gpio<13>
rlabel metal1 -110746 51273 -103746 58273 0 gpio<14>
rlabel metal1 168188 302860 175188 309860 0 adc1_in
rlabel metal1 151388 302860 158388 309860 0 adc0_in
rlabel metal1 247838 71885 254838 78885 0 comp_inp
rlabel metal1 247838 88685 254838 95685 0 comp_inn
rlabel space 185022 302827 192022 309827 0 adc_low
rlabel space 201822 302827 208822 309827 0 adc_high
rlabel space 218622 302827 225622 309827 0 analog_out
<< end >>
