magic
tech EFXH018D
magscale 1 2
timestamp 1567010579
<< error_s >>
rect -94573 327167 -94173 333967
rect -77773 327167 -77373 333967
rect -60973 327167 -60573 333967
rect -44173 327167 -43773 333967
rect -27373 327167 -26973 333967
rect -10573 327167 -10173 333967
rect 6227 327167 6627 333967
rect 23027 327167 23427 333967
rect 33027 327167 33427 333967
rect 43027 327167 43427 333967
rect 53027 327167 53427 333967
rect 63027 327167 63427 333967
rect 79827 327167 80227 333967
rect 96627 327167 97027 333967
rect 106627 327167 107027 333967
rect 123427 327167 123827 333967
rect 140227 327167 140627 333967
rect 157027 327167 157427 333967
rect 167027 327167 167427 333967
rect 177027 327167 177427 333967
rect 187027 327167 187427 333967
rect 197027 327167 197427 333967
rect 206927 327167 207427 333967
rect 299627 327167 300127 333967
rect 316427 327167 316827 333967
rect 333227 327167 333627 333967
rect 337227 327167 337627 333967
rect 339227 327167 339627 333967
rect 356027 327167 356427 333967
rect 217829 322654 222353 322682
rect 217829 316311 217857 322654
rect 222325 316311 222353 322654
rect 217829 316283 222353 316311
rect 284101 322386 288491 322414
rect 284101 316311 284129 322386
rect 288463 316311 288491 322386
rect 284101 316283 288491 316311
rect -94573 305543 -94173 311943
rect -77773 305543 -77373 311943
rect -60973 305543 -60573 311943
rect -44173 305543 -43773 311943
rect -27373 305543 -26973 311943
rect -10573 305543 -10173 311943
rect 6227 305543 6627 311943
rect 23027 305543 23427 311943
rect 33027 305543 33427 311943
rect 43027 305543 43427 311943
rect 53027 305543 53427 311943
rect 63027 305543 63427 311943
rect 79827 305543 80227 311943
rect 96627 305543 97027 311943
rect 106627 305543 107027 311943
rect 123427 305543 123827 311943
rect 140227 305543 140627 311943
rect 157027 305543 157427 311943
rect 167027 305543 167427 311943
rect 177027 305543 177427 311943
rect 187027 305543 187427 311943
rect 197027 305543 197427 311943
rect 206927 305543 207427 311943
rect 299627 305543 300127 311943
rect 316427 305543 316827 311943
rect 333227 305543 333627 311943
rect 337227 305543 337627 311943
rect 339227 305543 339627 311943
rect 356027 305543 356427 311943
rect -94773 304315 -94173 305043
rect -77973 304315 -77373 305043
rect -61173 304315 -60573 305043
rect -44373 304315 -43773 305043
rect -27573 304315 -26973 305043
rect -10773 304315 -10173 305043
rect 6027 304315 6627 305043
rect 22827 304315 23427 305043
rect 32827 304315 33427 305043
rect 42827 304315 43427 305043
rect 52827 304315 53427 305043
rect 62827 304315 63427 305043
rect 79627 304315 80227 305043
rect 96427 304315 97027 305043
rect 106427 304315 107027 305043
rect 123227 304315 123827 305043
rect 140027 304315 140627 305043
rect 156827 304315 157427 305043
rect 166827 304315 167427 305043
rect 176827 304315 177427 305043
rect 186827 304315 187427 305043
rect 196827 304315 197427 305043
rect 206827 304315 207427 305043
rect 299527 304315 300127 305043
rect 316227 304315 316827 305043
rect 333027 304315 333627 305043
rect 337027 304315 337627 305043
rect 339027 304315 339627 305043
rect 355827 304315 356427 305043
rect -94773 303215 -94173 303815
rect -77973 303215 -77373 303815
rect -61173 303215 -60573 303815
rect -44373 303215 -43773 303815
rect -27573 303215 -26973 303815
rect -10773 303215 -10173 303815
rect 6027 303215 6627 303815
rect 22827 303215 23427 303815
rect 32827 303215 33427 303815
rect 42827 303215 43427 303815
rect 52827 303215 53427 303815
rect 62827 303215 63427 303815
rect 79627 303215 80227 303815
rect 96427 303215 97027 303815
rect 106427 303215 107027 303815
rect 123227 303215 123827 303815
rect 140027 303215 140627 303815
rect 156827 303215 157427 303815
rect 166827 303215 167427 303815
rect 176827 303215 177427 303815
rect 186827 303215 187427 303815
rect 196827 303215 197427 303815
rect 206827 303215 207427 303815
rect 299527 303215 300127 303815
rect 316227 303215 316827 303815
rect 333027 303215 333627 303815
rect 337027 303215 337627 303815
rect 339027 303215 339627 303815
rect 355827 303215 356427 303815
rect -126673 302067 -119873 302467
rect -104649 302067 -98249 302467
rect -97749 301867 -97021 302467
rect -96521 301867 -95921 302467
rect -95421 301867 -94821 302467
rect -94773 302115 -94173 302715
rect -77973 302115 -77373 302715
rect -61173 302115 -60573 302715
rect -44373 302115 -43773 302715
rect -27573 302115 -26973 302715
rect -10773 302115 -10173 302715
rect 6027 302115 6627 302715
rect 22827 302115 23427 302715
rect 32827 302115 33427 302715
rect 42827 302115 43427 302715
rect 52827 302115 53427 302715
rect 62827 302115 63427 302715
rect 79627 302115 80227 302715
rect 96427 302115 97027 302715
rect 106427 302115 107027 302715
rect 123227 302115 123827 302715
rect 140027 302115 140627 302715
rect 156827 302115 157427 302715
rect 166827 302115 167427 302715
rect 176827 302115 177427 302715
rect 186827 302115 187427 302715
rect 196827 302115 197427 302715
rect 206827 302115 207427 302715
rect 299527 302115 300127 302715
rect 316227 302115 316827 302715
rect 333027 302115 333627 302715
rect 337027 302115 337627 302715
rect 339027 302115 339627 302715
rect 355827 302467 356427 302715
rect 355827 302115 356675 302467
rect 356075 301867 356675 302115
rect 357175 301867 357775 302467
rect 358275 301867 359003 302467
rect 359503 302067 365903 302467
rect 381127 302067 387927 302467
rect -126673 285267 -119873 285667
rect -104649 285267 -98249 285667
rect -97749 285067 -97021 285667
rect -96521 285067 -95921 285667
rect -95421 285067 -94821 285667
rect 356075 285067 356675 285667
rect 357175 285067 357775 285667
rect 358275 285067 359003 285667
rect 359503 285267 365903 285667
rect 381127 285267 387927 285667
rect -126673 268467 -119873 268867
rect -104649 268467 -98249 268867
rect -97749 268267 -97021 268867
rect -96521 268267 -95921 268867
rect -95421 268267 -94821 268867
rect 356075 268267 356675 268867
rect 357175 268267 357775 268867
rect 358275 268267 359003 268867
rect 359503 268467 365903 268867
rect 381127 268467 387927 268867
rect -126673 258467 -119873 258867
rect -104649 258467 -98249 258867
rect -97749 258267 -97021 258867
rect -96521 258267 -95921 258867
rect -95421 258267 -94821 258867
rect 356075 251467 356675 252067
rect 357175 251467 357775 252067
rect 358275 251467 359003 252067
rect 359503 251667 365903 252067
rect 381127 251667 387927 252067
rect -126673 241667 -119873 242067
rect -104649 241667 -98249 242067
rect -97749 241467 -97021 242067
rect -96521 241467 -95921 242067
rect -95421 241467 -94821 242067
rect 356075 234667 356675 235267
rect 357175 234667 357775 235267
rect 358275 234667 359003 235267
rect 359503 234867 365903 235267
rect 381127 234867 387927 235267
rect -126673 224867 -119873 225267
rect -104649 224867 -98249 225267
rect -97749 224667 -97021 225267
rect -96521 224667 -95921 225267
rect -95421 224667 -94821 225267
rect 356075 217867 356675 218467
rect 357175 217867 357775 218467
rect 358275 217867 359003 218467
rect 359503 218067 365903 218467
rect 381127 218067 387927 218467
rect -126673 208067 -119873 208467
rect -104649 208067 -98249 208467
rect -97749 207867 -97021 208467
rect -96521 207867 -95921 208467
rect -95421 207867 -94821 208467
rect 356075 207867 356675 208467
rect 357175 207867 357775 208467
rect 358275 207867 359003 208467
rect 359503 208067 365903 208467
rect 381127 208067 387927 208467
rect 356075 197867 356675 198467
rect 357175 197867 357775 198467
rect 358275 197867 359003 198467
rect 359503 198067 365903 198467
rect 381127 198067 387927 198467
rect -126673 191267 -119873 191667
rect -104649 191267 -98249 191667
rect -97749 191067 -97021 191667
rect -96521 191067 -95921 191667
rect -95421 191067 -94821 191667
rect 356075 187867 356675 188467
rect 357175 187867 357775 188467
rect 358275 187867 359003 188467
rect 359503 188067 365903 188467
rect 381127 188067 387927 188467
rect -96521 180667 -95921 181267
rect -95421 180667 -94821 181267
rect -126673 178867 -119873 179267
rect -104649 178867 -98249 179267
rect -97749 178667 -97021 179267
rect -96521 178667 -95921 179267
rect -95421 178667 -94821 179267
rect 356075 177867 356675 178467
rect 357175 177867 357775 178467
rect 358275 177867 359003 178467
rect 359503 178067 365903 178467
rect 381127 178067 387927 178467
rect -126673 162067 -119873 162467
rect -104649 162067 -98249 162467
rect -97749 161867 -97021 162467
rect -96521 161867 -95921 162467
rect -95421 161867 -94821 162467
rect 356075 161067 356675 161667
rect 357175 161067 357775 161667
rect 358275 161067 359003 161667
rect 359503 161267 365903 161667
rect 381127 161267 387927 161667
rect -126673 145267 -119873 145667
rect -104649 145267 -98249 145667
rect -97749 145067 -97021 145667
rect -96521 145067 -95921 145667
rect -95421 145067 -94821 145667
rect 356075 144267 356675 144867
rect 357175 144267 357775 144867
rect 358275 144267 359003 144867
rect 359503 144467 365903 144867
rect 381127 144467 387927 144867
rect 356075 134267 356675 134867
rect 357175 134267 357775 134867
rect 358275 134267 359003 134867
rect 359503 134467 365903 134867
rect 381127 134467 387927 134867
rect -126673 128467 -119873 128867
rect -104649 128467 -98249 128867
rect -97749 128267 -97021 128867
rect -96521 128267 -95921 128867
rect -95421 128267 -94821 128867
rect 356075 117467 356675 118067
rect 357175 117467 357775 118067
rect 358275 117467 359003 118067
rect 359503 117667 365903 118067
rect 381127 117667 387927 118067
rect -126673 111667 -119873 112067
rect -104649 111667 -98249 112067
rect -97749 111467 -97021 112067
rect -96521 111467 -95921 112067
rect -95421 111467 -94821 112067
rect 356075 100667 356675 101267
rect 357175 100667 357775 101267
rect 358275 100667 359003 101267
rect 359503 100867 365903 101267
rect 381127 100867 387927 101267
rect -126673 94867 -119873 95267
rect -104649 94867 -98249 95267
rect -97749 94667 -97021 95267
rect -96521 94667 -95921 95267
rect -95421 94667 -94821 95267
rect 356075 90667 356675 91267
rect 357175 90667 357775 91267
rect 358275 90667 359003 91267
rect 359503 90867 365903 91267
rect 381127 90867 387927 91267
rect 356075 80667 356675 81267
rect 357175 80667 357775 81267
rect 358275 80667 359003 81267
rect 359503 80867 365903 81267
rect 381127 80867 387927 81267
rect -126673 78067 -119873 78467
rect -104649 78067 -98249 78467
rect -97749 77867 -97021 78467
rect -96521 77867 -95921 78467
rect -95421 77867 -94821 78467
rect 356075 70667 356675 71267
rect 357175 70667 357775 71267
rect 358275 70667 359003 71267
rect 359503 70867 365903 71267
rect 381127 70867 387927 71267
rect -126673 61267 -119873 61667
rect -104649 61267 -98249 61667
rect -97749 61067 -97021 61667
rect -96521 61067 -95921 61667
rect -95421 61067 -94821 61667
rect 356075 53867 356675 54467
rect 357175 53867 357775 54467
rect 358275 53867 359003 54467
rect 359503 54067 365903 54467
rect 381127 54067 387927 54467
rect -126673 51267 -119873 51667
rect -104649 51267 -98249 51667
rect -97749 51067 -97021 51667
rect -96521 51067 -95921 51667
rect -95421 51067 -94821 51667
rect 356075 37067 356675 37667
rect 357175 37067 357775 37667
rect 358275 37067 359003 37667
rect 359503 37267 365903 37667
rect 381127 37267 387927 37667
rect -126673 34467 -119873 34967
rect -104649 34467 -98249 34967
rect -97749 34367 -97021 34967
rect -96521 34367 -95921 34967
rect -95421 34367 -94821 34967
rect -114102 27699 -110225 27727
rect -114102 24415 -114074 27699
rect -110253 24415 -110225 27699
rect 356075 27067 356675 27667
rect 357175 27067 357775 27667
rect 358275 27067 359003 27667
rect 359503 27267 365903 27667
rect 381127 27267 387927 27667
rect -114102 24387 -110225 24415
rect 356075 17067 356675 17667
rect 357175 17067 357775 17667
rect 358275 17067 359003 17667
rect 359503 17267 365903 17667
rect 381127 17267 387927 17667
rect 356075 7067 356675 7667
rect 357175 7067 357775 7667
rect 358275 7067 359003 7667
rect 359503 7267 365903 7667
rect 381127 7267 387927 7667
rect 356075 -2933 356675 -2333
rect 357175 -2933 357775 -2333
rect 358275 -2933 359003 -2333
rect 359503 -2733 365903 -2333
rect 381127 -2733 387927 -2333
rect -114520 -10941 -110046 -10913
rect -114520 -14465 -114492 -10941
rect -110074 -14465 -110046 -10941
rect -114520 -14493 -110046 -14465
rect 356075 -19733 356675 -19133
rect 357175 -19733 357775 -19133
rect 358275 -19733 359003 -19133
rect 359503 -19533 365903 -19133
rect 381127 -19533 387927 -19133
rect -98673 -20333 -94791 -20133
rect -126673 -20833 -119873 -20333
rect -104649 -20541 -94791 -20333
rect -104649 -20833 -98249 -20541
rect -98157 -20833 -97996 -20541
rect -97904 -20833 -96660 -20541
rect -96540 -20633 -95620 -20541
rect -95501 -20633 -94821 -20541
rect -96540 -20833 -94821 -20633
rect -98673 -20933 -98249 -20833
rect -97749 -20933 -97021 -20833
rect -96521 -20933 -95921 -20833
rect -95421 -20933 -94821 -20833
rect 356075 -36533 356675 -35933
rect 357175 -36533 357775 -35933
rect 358275 -36533 359003 -35933
rect 359503 -36333 365903 -35933
rect 381127 -36333 387927 -35933
rect -126673 -37533 -119873 -37133
rect -104649 -37533 -98249 -37133
rect -97749 -37733 -97021 -37133
rect -96521 -37733 -95921 -37133
rect -95421 -37733 -94821 -37133
rect 356075 -46733 356675 -46133
rect 357175 -46733 357775 -46133
rect 358275 -46733 359003 -46133
rect 359503 -46333 365903 -46133
rect 381127 -46333 387927 -46133
rect -126673 -47533 -119873 -47133
rect -104649 -47533 -98249 -47133
rect -97749 -47733 -97021 -47133
rect -96521 -47733 -95921 -47133
rect -95421 -47733 -94821 -47133
rect -7673 -47689 -7073 -47476
rect -7481 -47781 -7073 -47689
rect -94773 -48381 -94173 -47781
rect -93773 -48381 -93173 -47781
rect -92673 -48381 -92073 -47781
rect -75973 -48381 -75373 -47781
rect -59173 -48381 -58573 -47781
rect -42373 -48381 -41773 -47781
rect -25573 -48381 -24973 -47781
rect -8773 -48381 -8173 -47781
rect -7673 -48461 -7073 -47781
rect -7673 -48580 -7573 -48461
rect -7481 -48580 -7073 -48461
rect -94773 -49481 -94173 -48881
rect -93773 -49481 -93173 -48881
rect -92673 -49481 -92073 -48881
rect -75973 -49481 -75373 -48881
rect -59173 -49481 -58573 -48881
rect -42373 -49481 -41773 -48881
rect -25573 -49481 -24973 -48881
rect -8773 -49481 -8173 -48881
rect -7673 -48980 -7073 -48580
rect -7673 -49100 -7573 -48980
rect -7481 -49100 -7073 -48980
rect -7673 -49500 -7073 -49100
rect -7481 -49620 -7073 -49500
rect -94773 -50709 -94173 -49981
rect -93773 -50709 -93173 -49981
rect -92673 -50709 -92073 -49981
rect -75973 -50709 -75373 -49981
rect -59173 -50709 -58573 -49981
rect -42373 -50709 -41773 -49981
rect -25573 -50709 -24973 -49981
rect -8773 -50709 -8173 -49981
rect -7673 -50300 -7073 -49620
rect -7673 -50392 -7573 -50300
rect -7481 -50392 -7073 -50300
rect -7673 -50576 -7073 -50392
rect -7673 -50668 -7573 -50576
rect -7481 -50668 -7073 -50576
rect -7673 -50864 -7073 -50668
rect -7481 -50956 -7073 -50864
rect -7673 -51117 -7073 -50956
rect -7481 -51209 -7073 -51117
rect -94573 -57609 -94173 -51209
rect -93673 -57609 -93173 -51209
rect -92573 -57609 -92073 -51209
rect -75773 -57609 -75373 -51209
rect -58973 -57609 -58573 -51209
rect -42173 -57609 -41773 -51209
rect -25373 -57609 -24973 -51209
rect -8673 -57609 -8173 -51209
rect -7673 -57609 -7073 -51209
rect -7481 -57701 -7073 -57609
rect -7673 -58109 -7073 -57701
rect 84327 -47689 84927 -47476
rect 84327 -47781 84735 -47689
rect 356075 -47733 356675 -47133
rect 357175 -47733 357775 -47133
rect 358275 -47733 359003 -47133
rect 359503 -47533 365903 -47133
rect 381127 -47533 387927 -47133
rect 84327 -48381 85427 -47781
rect 92827 -48381 93427 -47781
rect 93827 -48381 94427 -47781
rect 103827 -48381 104427 -47781
rect 120627 -48381 121227 -47781
rect 130627 -48381 131227 -47781
rect 140627 -48381 141227 -47781
rect 157427 -48381 158027 -47781
rect 174227 -48381 174827 -47781
rect 184227 -48381 184827 -47781
rect 201027 -48381 201627 -47781
rect 217827 -48381 218427 -47781
rect 227827 -48381 228427 -47781
rect 237827 -48381 238427 -47781
rect 254627 -48381 255227 -47781
rect 271427 -48381 272027 -47781
rect 288227 -48381 288827 -47781
rect 305027 -48381 305627 -47781
rect 321827 -48381 322427 -47781
rect 331827 -48381 332427 -47781
rect 335827 -48381 336427 -47781
rect 337827 -48381 338427 -47781
rect 338827 -48381 339427 -47781
rect 355827 -48381 356427 -47781
rect 84327 -48881 84735 -48381
rect 84827 -48881 85527 -48381
rect 84327 -49100 85527 -48881
rect 84327 -49481 85427 -49100
rect 92827 -49481 93427 -48881
rect 93827 -49481 94427 -48881
rect 103827 -49481 104427 -48881
rect 120627 -49481 121227 -48881
rect 130627 -49481 131227 -48881
rect 140627 -49481 141227 -48881
rect 157427 -49481 158027 -48881
rect 174227 -49481 174827 -48881
rect 184227 -49481 184827 -48881
rect 201027 -49481 201627 -48881
rect 217827 -49481 218427 -48881
rect 227827 -49481 228427 -48881
rect 237827 -49481 238427 -48881
rect 254627 -49481 255227 -48881
rect 271427 -49481 272027 -48881
rect 288227 -49481 288827 -48881
rect 305027 -49481 305627 -48881
rect 321827 -49481 322427 -48881
rect 331827 -49481 332427 -48881
rect 335827 -49481 336427 -48881
rect 337827 -49481 338427 -48881
rect 338827 -49481 339427 -48881
rect 355827 -49481 356427 -48881
rect 84327 -50109 84735 -49481
rect 84827 -49500 85427 -49481
rect 84827 -49700 85427 -49620
rect 84827 -50109 85527 -49700
rect 84327 -50668 85527 -50109
rect 84327 -50709 85427 -50668
rect 92827 -50709 93427 -49981
rect 93827 -50709 94427 -49981
rect 103827 -50709 104427 -49981
rect 120627 -50709 121227 -49981
rect 130627 -50709 131227 -49981
rect 140627 -50709 141227 -49981
rect 157427 -50709 158027 -49981
rect 174227 -50709 174827 -49981
rect 184227 -50709 184827 -49981
rect 201027 -50709 201627 -49981
rect 217827 -50709 218427 -49981
rect 227827 -50709 228427 -49981
rect 237827 -50709 238427 -49981
rect 254627 -50709 255227 -49981
rect 271427 -50709 272027 -49981
rect 288227 -50709 288827 -49981
rect 305027 -50709 305627 -49981
rect 321827 -50709 322427 -49981
rect 331827 -50709 332427 -49981
rect 335827 -50709 336427 -49981
rect 337827 -50709 338427 -49981
rect 338827 -50709 339427 -49981
rect 355827 -50709 356427 -49981
rect 84327 -50956 84735 -50709
rect 84827 -50864 85427 -50709
rect 84327 -51117 84927 -50956
rect 84327 -57701 84735 -51117
rect 84827 -57609 85427 -51209
rect 93027 -57609 93427 -51209
rect 94027 -57609 94427 -51209
rect 104027 -57609 104427 -51209
rect 120827 -57609 121227 -51209
rect 130827 -57609 131227 -51209
rect 140827 -57609 141227 -51209
rect 157627 -57609 158027 -51209
rect 174427 -57609 174827 -51209
rect 184427 -57609 184827 -51209
rect 201227 -57609 201627 -51209
rect 218027 -57609 218427 -51209
rect 228027 -57609 228427 -51209
rect 238027 -57609 238427 -51209
rect 254827 -57609 255227 -51209
rect 271627 -57609 272027 -51209
rect 288427 -57609 288827 -51209
rect 305227 -57609 305627 -51209
rect 322027 -57609 322427 -51209
rect 332027 -57609 332427 -51209
rect 336027 -57609 336427 -51209
rect 338027 -57609 338427 -51209
rect 339227 -57609 339427 -51209
rect 356027 -57609 356427 -51209
rect 84327 -58109 84927 -57701
rect 2983 -61977 8133 -61569
rect 2983 -68052 3391 -61977
rect 3483 -62477 7633 -62069
rect 3483 -67552 3891 -62477
rect 7225 -67552 7633 -62477
rect 3483 -67960 7633 -67552
rect 7725 -68052 8133 -61977
rect 2983 -68460 8133 -68052
rect 69121 -61977 74405 -61569
rect 69121 -68320 69529 -61977
rect 69621 -62477 73905 -62069
rect 69621 -67820 70029 -62477
rect 73497 -67820 73905 -62477
rect 69621 -68228 73905 -67820
rect 73997 -68320 74405 -61977
rect 69121 -68728 74405 -68320
rect -7673 -72741 -7073 -72333
rect -7481 -72833 -7073 -72741
rect -94573 -79633 -94173 -72833
rect -93673 -79633 -93173 -72833
rect -92573 -79633 -92073 -72833
rect -75773 -79633 -75373 -72833
rect -58973 -79633 -58573 -72833
rect -42173 -79633 -41773 -72833
rect -25373 -79633 -24973 -72833
rect -8673 -79633 -8173 -72833
rect -7673 -79633 -7073 -72833
rect 84327 -72741 84927 -72333
rect 84327 -79633 84735 -72741
rect 84827 -79633 85427 -72833
rect 93027 -79633 93427 -72833
rect 94027 -79633 94427 -72833
rect 104027 -79633 104427 -72833
rect 120827 -79633 121227 -72833
rect 130827 -79633 131227 -72833
rect 140827 -79633 141227 -72833
rect 157627 -79633 158027 -72833
rect 174427 -79633 174827 -72833
rect 184427 -79633 184827 -72833
rect 201227 -79633 201627 -72833
rect 218027 -79633 218427 -72833
rect 228027 -79633 228427 -72833
rect 238027 -79633 238427 -72833
rect 254827 -79633 255227 -72833
rect 271627 -79633 272027 -72833
rect 288427 -79633 288827 -72833
rect 305227 -79633 305627 -72833
rect 322027 -79633 322427 -72833
rect 332027 -79633 332427 -72833
rect 336027 -79633 336427 -72833
rect 338027 -79633 338427 -72833
rect 339227 -79633 339427 -72833
rect 356027 -79633 356427 -72833
<< metal1 >>
rect -89307 314732 -82676 323657
rect -73117 315671 -66660 323257
rect -56317 315671 -49860 323257
rect -39517 315671 -33060 323257
rect -22717 315671 -16260 323257
rect -5917 315671 540 323257
rect 10883 315671 17340 323257
rect 67929 315690 74386 323276
rect 84729 315690 91186 323276
rect 111529 315690 117986 323276
rect 128329 315690 134786 323276
rect 145129 315690 151586 323276
rect 218762 317000 221057 321592
rect 285132 317000 287427 321592
rect 304823 316062 310764 323116
rect 321623 316062 327564 323116
rect 344449 316120 350390 323174
rect -116217 290579 -108447 296323
rect 369053 289951 377601 296125
rect -117641 273192 -108233 279730
rect 369940 274803 376306 279297
rect 370002 256958 377759 262815
rect -117320 245880 -107876 253893
rect 369211 240020 378076 246035
rect -117455 229677 -107460 236387
rect 369053 223557 378234 229256
rect -117455 212877 -107460 219587
rect -117312 196029 -107603 203168
rect -117155 166595 -107704 173799
rect 369816 167810 376581 172461
rect -117310 149977 -107859 157181
rect 368979 149924 377408 155403
rect -116941 133772 -107241 140318
rect -116558 116854 -107853 123653
rect 368961 122718 377921 129374
rect 369393 106440 376581 111514
rect -117256 100525 -108391 105591
rect -116705 82589 -107714 89766
rect -116623 66966 -108391 72664
rect 368450 58703 377782 65962
rect -117397 39351 -107728 45931
rect 368450 41903 377782 49162
rect 369451 -13575 377901 -8217
rect -117178 -32710 -107083 -25770
rect 368504 -31678 377782 -24769
rect -87393 -69600 -81084 -60847
rect -70290 -69844 -63641 -61138
rect -54460 -69686 -46703 -60979
rect -37838 -69686 -30715 -61613
rect -20650 -69433 -14256 -60528
rect 4145 -67471 6518 -62988
rect 70472 -67471 72977 -62856
rect 108500 -70049 115641 -60687
rect 145300 -70049 152441 -60687
rect 162121 -70366 169420 -60369
rect 189047 -70078 196132 -60189
rect 205726 -70078 212811 -60779
rect 242746 -69468 249188 -61026
rect 259629 -69690 265850 -60803
rect 276513 -69912 282956 -60803
rect 293175 -69690 300062 -61026
rect 309697 -70150 316892 -60731
rect 344225 -69745 350147 -62244
<< metaltpl >>
rect -113603 24811 -110754 27289
rect -114081 -13937 -111232 -11459
use CORNERESDF  CORNERESDF_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -126673 -1 0 333967
box 0 0 32000 32000
use BBCUD4F  GPIO_buf_11 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform -1 0 -77873 0 -1 333967
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_10
timestamp 1529526440
transform -1 0 -61073 0 -1 333967
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_9
timestamp 1529526440
transform -1 0 -44273 0 -1 333967
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_8
timestamp 1529526440
transform -1 0 -27473 0 -1 333967
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_7
timestamp 1529526440
transform -1 0 -10673 0 -1 333967
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_6
timestamp 1529526440
transform -1 0 6127 0 -1 333967
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_5
timestamp 1529526440
transform -1 0 22927 0 -1 333967
box 0 0 16800 32000
use FILLER50F  FILLER50F_30 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform -1 0 32927 0 -1 333967
box 0 0 10000 32000
use FILLER50F  FILLER50F_23
timestamp 1529526440
transform -1 0 42927 0 -1 333967
box 0 0 10000 32000
use FILLER50F  FILLER50F_18
timestamp 1529526440
transform -1 0 52927 0 -1 333967
box 0 0 10000 32000
use FILLER50F  FILLER50F_19
timestamp 1529526440
transform -1 0 62927 0 -1 333967
box 0 0 10000 32000
use BBCUD4F  GPIO_buf_4
timestamp 1529526440
transform -1 0 79727 0 -1 333967
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_3
timestamp 1529526440
transform -1 0 96527 0 -1 333967
box 0 0 16800 32000
use FILLER50F  FILLER50F_20
timestamp 1529526440
transform -1 0 106527 0 -1 333967
box 0 0 10000 32000
use BBCUD4F  GPIO_buf_2
timestamp 1529526440
transform -1 0 123327 0 -1 333967
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_1
timestamp 1529526440
transform -1 0 140127 0 -1 333967
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_0
timestamp 1529526440
transform -1 0 156927 0 -1 333967
box 0 0 16800 32000
use FILLER50F  FILLER50F_15
timestamp 1529526440
transform -1 0 166927 0 -1 333967
box 0 0 10000 32000
use FILLER50F  FILLER50F_16
timestamp 1529526440
transform -1 0 176927 0 -1 333967
box 0 0 10000 32000
use FILLER50F  FILLER50F_17
timestamp 1529526440
transform -1 0 186927 0 -1 333967
box 0 0 10000 32000
use FILLER50F  FILLER50F_24
timestamp 1529526440
transform -1 0 196927 0 -1 333967
box 0 0 10000 32000
use FILLER50F  FILLER50F_25
timestamp 1529526440
transform -1 0 206927 0 -1 333967
box 0 0 10000 32000
use VDDORPADF  vddor_pad_3 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -126673 -1 0 301967
box 0 0 16800 32000
use GNDORPADF  gndor_pad_4 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -126673 -1 0 285167
box 0 0 16800 32000
use FILLER50F  FILLER50F_2
timestamp 1529526440
transform 0 1 -126673 -1 0 268367
box 0 0 10000 32000
use aregc01_3v3  regulator2 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1516677094
transform -1 0 299527 0 -1 333967
box 0 0 92600 70740
use VDDORPADF  vddor_pad_0
timestamp 1529526440
transform -1 0 316327 0 -1 333967
box 0 0 16800 32000
use GNDORPADF  gndor_pad_1
timestamp 1529526440
transform -1 0 333127 0 -1 333967
box 0 0 16800 32000
use FILLER20F  FILLER20F_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform -1 0 337127 0 -1 333967
box 0 0 4000 32000
use FILLER10F  FILLER10F_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform -1 0 339127 0 -1 333967
box 0 0 2000 32000
use VDDORPADF  vddor_pad_1
timestamp 1529526440
transform -1 0 355927 0 -1 333967
box 0 0 16800 32000
use CORNERESDF  CORNERESDF_0
timestamp 1529526440
transform -1 0 387927 0 -1 333967
box 0 0 32000 32000
use ICF  spi_master_sdi_buf /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 -1 387927 1 0 285167
box 0 0 16800 32000
use GNDORPADF  gndor_pad_2
timestamp 1529526440
transform 0 -1 387927 1 0 268367
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_12
timestamp 1529526440
transform 0 1 -126673 -1 0 258367
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_13
timestamp 1529526440
transform 0 1 -126673 -1 0 241567
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_14
timestamp 1529526440
transform 0 1 -126673 -1 0 224767
box 0 0 16800 32000
use BBCUD4F  GPIO_buf_15
timestamp 1529526440
transform 0 1 -126673 -1 0 207967
box 0 0 16800 32000
use FILLER50F  FILLER50F_22
timestamp 1529526440
transform 0 1 -126673 -1 0 191167
box 0 0 10000 32000
use FILLER02F  FILLER02F_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -126673 -1 0 181167
box 0 0 400 32000
use FILLER10F  FILLER10F_1
timestamp 1529526440
transform 0 1 -126673 -1 0 180767
box 0 0 2000 32000
use APR00DF  comp_inp_pad /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 1 -126673 -1 0 178767
box 0 0 16800 32000
use APR00DF  comp_inn_pad
timestamp 1529526440
transform 0 1 -126673 -1 0 161967
box 0 0 16800 32000
use APR00DF  ana_out_pad
timestamp 1529526440
transform 0 1 -126673 -1 0 145167
box 0 0 16800 32000
use APR00DF  adc_high_pad
timestamp 1529526440
transform 0 1 -126673 -1 0 128367
box 0 0 16800 32000
use APR00DF  adc_low_pad
timestamp 1529526440
transform 0 1 -126673 -1 0 111567
box 0 0 16800 32000
use APR00DF  adc1_pad
timestamp 1529526440
transform 0 1 -126673 -1 0 94767
box 0 0 16800 32000
use APR00DF  adc0_pad
timestamp 1529526440
transform 0 1 -126673 -1 0 77967
box 0 0 16800 32000
use FILLER50F  FILLER50F_21
timestamp 1529526440
transform 0 1 -126673 -1 0 61167
box 0 0 10000 32000
use APR00DF  nvref_ext_pad
timestamp 1529526440
transform 0 1 -126673 -1 0 51167
box 0 0 16800 32000
use BT4F  spi_master_csb_buf /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 -1 387927 1 0 251567
box 0 0 16800 32000
use BT4F  spi_master_sck_buf
timestamp 1529526440
transform 0 -1 387927 1 0 234767
box 0 0 16800 32000
use BT4F  spi_master_sdo_buf
timestamp 1529526440
transform 0 -1 387927 1 0 217967
box 0 0 16800 32000
use FILLER50F  FILLER50F_31
timestamp 1529526440
transform 0 -1 387927 1 0 207967
box 0 0 10000 32000
use FILLER50F  FILLER50F_14
timestamp 1529526440
transform 0 -1 387927 1 0 197967
box 0 0 10000 32000
use FILLER50F  FILLER50F_13
timestamp 1529526440
transform 0 -1 387927 1 0 187967
box 0 0 10000 32000
use FILLER50F  FILLER50F_12
timestamp 1529526440
transform 0 -1 387927 1 0 177967
box 0 0 10000 32000
use ICF  ser_rx_buf
timestamp 1529526440
transform 0 -1 387927 1 0 161167
box 0 0 16800 32000
use BT4F  ser_tx_buf
timestamp 1529526440
transform 0 -1 387927 1 0 144367
box 0 0 16800 32000
use FILLER50F  FILLER50F_33
timestamp 1529526440
transform 0 -1 387927 1 0 134367
box 0 0 10000 32000
use VDDPADF  vdd_pad_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 -1 387927 1 0 117567
box 0 0 16800 32000
use GNDORPADF  gndor_pad_0
timestamp 1529526440
transform 0 -1 387927 1 0 100767
box 0 0 16800 32000
use FILLER50F  FILLER50F_6
timestamp 1529526440
transform 0 -1 387927 1 0 90767
box 0 0 10000 32000
use FILLER50F  FILLER50F_5
timestamp 1529526440
transform 0 -1 387927 1 0 80767
box 0 0 10000 32000
use FILLER50F  FILLER50F_1
timestamp 1529526440
transform 0 -1 387927 1 0 70767
box 0 0 10000 32000
use BBCUD4F  i2c_scl_pad
timestamp 1529526440
transform 0 -1 387927 1 0 53967
box 0 0 16800 32000
use BBCUD4F  i2c_sda_pad
timestamp 1529526440
transform 0 -1 387927 1 0 37167
box 0 0 16800 32000
use axtoc02_3v3  xtal /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/A_CELLS_3V3
timestamp 1516677002
transform 0 1 -126673 -1 0 34367
box 0 0 55200 31882
use FILLER50F  FILLER50F_36
timestamp 1529526440
transform 0 -1 387927 1 0 27167
box 0 0 10000 32000
use FILLER50F  FILLER50F_37
timestamp 1529526440
transform 0 -1 387927 1 0 17167
box 0 0 10000 32000
use FILLER50F  FILLER50F_38
timestamp 1529526440
transform 0 -1 387927 1 0 7167
box 0 0 10000 32000
use FILLER50F  FILLER50F_39
timestamp 1529526440
transform 0 -1 387927 1 0 -2833
box 0 0 10000 32000
use VDDORPADF  vddor_pad_2
timestamp 1529526440
transform 0 1 -126673 -1 0 -20833
box 0 0 16800 32000
use FILLER50F  FILLER50F_7
timestamp 1529526440
transform 0 1 -126673 -1 0 -37633
box 0 0 10000 32000
use CORNERESDF  CORNERESDF_2
timestamp 1529526440
transform 1 0 -126673 0 1 -79633
box 0 0 32000 32000
use FILLER05F  FILLER05F_3 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 1 0 -94673 0 1 -79633
box 0 0 1000 32000
use POWERCUTVDD3FC  pwr_cut_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_FC3V
timestamp 1516645956
transform -1 0 -92673 0 1 -79633
box 0 0 1000 32000
use BT4FC  sdo_buf /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_FC3V
timestamp 1529532354
transform 1 0 -92673 0 1 -79633
box 0 0 16800 32000
use ICFC  sdi_buf /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_FC3V
timestamp 1529532354
transform 1 0 -75873 0 1 -79633
box 0 0 16800 32000
use ICFC  csb_buf
timestamp 1529532354
transform 1 0 -59073 0 1 -79633
box 0 0 16800 32000
use ICFC  sck_buf
timestamp 1529532354
transform 1 0 -42273 0 1 -79633
box 0 0 16800 32000
use VDDPADFC  vdd3_pad /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_FC3V
timestamp 1529532354
transform 1 0 -25473 0 1 -79633
box 0 0 16800 32000
use POWERCUTVDD3FC  pwr_cut_1
timestamp 1516645956
transform 1 0 -8673 0 1 -79633
box 0 0 1000 32000
use aregc01_3v3  regulator1
timestamp 1516677094
transform 1 0 -7673 0 1 -79633
box 0 0 92600 70740
use GNDORPADF  GNDORPADF_1
timestamp 1529526440
transform 0 -1 387927 1 0 -19633
box 0 0 16800 32000
use ICF  irq_buf
timestamp 1529526440
transform 0 -1 387927 1 0 -36433
box 0 0 16800 32000
use FILLER50F  FILLER50F_40
timestamp 1529526440
transform 0 -1 387927 1 0 -46433
box 0 0 10000 32000
use FILLER01F  FILLER01F_1 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 0 -1 387927 1 0 -46633
box 0 0 200 32000
use FILLER05F  FILLER05F_1
timestamp 1529526440
transform 0 -1 387927 1 0 -47633
box 0 0 1000 32000
use FILLER40F  FILLER40F_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 1 0 84927 0 1 -79633
box 0 0 8000 32000
use FILLER05F  FILLER05F_2
timestamp 1529526440
transform 1 0 92927 0 1 -79633
box 0 0 1000 32000
use FILLER50F  FILLER50F_26
timestamp 1529526440
transform 1 0 93927 0 1 -79633
box 0 0 10000 32000
use GNDORPADF  gndor_pad_5
timestamp 1529526440
transform 1 0 103927 0 1 -79633
box 0 0 16800 32000
use FILLER50F  FILLER50F_32
timestamp 1529526440
transform 1 0 120727 0 1 -79633
box 0 0 10000 32000
use FILLER50F  FILLER50F_27
timestamp 1529526440
transform 1 0 130727 0 1 -79633
box 0 0 10000 32000
use VDDORPADF  vddor_pad_4
timestamp 1529526440
transform 1 0 140727 0 1 -79633
box 0 0 16800 32000
use VDDPADF  vdd_pad_1
timestamp 1529526440
transform 1 0 157527 0 1 -79633
box 0 0 16800 32000
use FILLER50F  FILLER50F_8
timestamp 1529526440
transform 1 0 174327 0 1 -79633
box 0 0 10000 32000
use BT4F  flash_clk_buf
timestamp 1529526440
transform 1 0 184327 0 1 -79633
box 0 0 16800 32000
use BT4F  flash_csb_buf
timestamp 1529526440
transform 1 0 201127 0 1 -79633
box 0 0 16800 32000
use FILLER50F  FILLER50F_28
timestamp 1529526440
transform 1 0 217927 0 1 -79633
box 0 0 10000 32000
use FILLER50F  FILLER50F_29
timestamp 1529526440
transform 1 0 227927 0 1 -79633
box 0 0 10000 32000
use BBC4F  flash_io_buf_0 /ef/tech/XFAB.3/EFXH018D/libs.ref/maglef/IO_CELLS_F3V
timestamp 1529526440
transform 1 0 237927 0 1 -79633
box 0 0 16800 32000
use BBC4F  flash_io_buf_1
timestamp 1529526440
transform 1 0 254727 0 1 -79633
box 0 0 16800 32000
use BBC4F  flash_io_buf_2
timestamp 1529526440
transform 1 0 271527 0 1 -79633
box 0 0 16800 32000
use BBC4F  flash_io_buf_3
timestamp 1529526440
transform 1 0 288327 0 1 -79633
box 0 0 16800 32000
use GNDORPADF  gndor_pad_3
timestamp 1529526440
transform 1 0 305127 0 1 -79633
box 0 0 16800 32000
use FILLER50F  FILLER50F_34
timestamp 1529526440
transform 1 0 321927 0 1 -79633
box 0 0 10000 32000
use FILLER20F  FILLER20F_1
timestamp 1529526440
transform 1 0 331927 0 1 -79633
box 0 0 4000 32000
use FILLER10F  FILLER10F_2
timestamp 1529526440
transform 1 0 335927 0 1 -79633
box 0 0 2000 32000
use FILLER05F  FILLER05F_0
timestamp 1529526440
transform 1 0 337927 0 1 -79633
box 0 0 1000 32000
use FILLER01F  FILLER01F_0
timestamp 1529526440
transform 1 0 338927 0 1 -79633
box 0 0 200 32000
use ICF  clk_ext_buf
timestamp 1529526440
transform 1 0 339127 0 1 -79633
box 0 0 16800 32000
use CORNERESDF  CORNERESDF_3
timestamp 1529526440
transform 0 -1 387927 1 0 -79633
box 0 0 32000 32000
<< labels >>
rlabel metal1 s 293175 -69690 300062 -61026 0 flash_io3
rlabel metal1 s 276513 -69912 282956 -60803 0 flash_io2
rlabel metal1 s 259629 -69690 265850 -60803 0 flash_io1
rlabel metal1 s 242746 -69468 249188 -61026 0 flash_io0
rlabel metal1 s 309697 -70150 316892 -60731 0 VSS
rlabel metal1 s 344225 -69745 350147 -62244 0 XCLK
rlabel metal1 s -117397 39351 -107728 45931 0 nvref_ext
rlabel metal1 s -117256 100525 -108391 105591 0 adc_low
rlabel metal1 s -116558 116854 -107853 123653 0 adc_high
rlabel metal1 s -117310 149977 -107859 157181 0 comp_inn
rlabel metal1 s -117155 166595 -107704 173799 0 comp_inp
rlabel metaltpl -114081 -13937 -111232 -11459 0 XO
rlabel metaltpl -113603 24811 -110754 27289 0 XI
rlabel metal1 s -116623 66966 -108391 72664 0 adc0_in
rlabel metal1 s -116941 133772 -107241 140318 0 analog_out
rlabel metal1 s -116705 82589 -107714 89766 0 adc1_in
rlabel metal1 -117178 -32710 -107083 -25770 0 VDD3V3
rlabel metal1 s 108500 -70049 115641 -60687 0 VSS
rlabel metal1 s 145300 -70049 152441 -60687 0 VDD3V3
rlabel metal1 s 162121 -70366 169420 -60369 0 VDD1V8
rlabel metal1 s 205726 -70078 212811 -60779 0 flash_csb
rlabel metal1 s 189047 -70078 196132 -60189 0 flash_clk
rlabel metal1 s 368450 41903 377782 49162 0 i2c_sda
rlabel metal1 s 368450 58703 377782 65962 0 i2c_scl
rlabel metal1 s 368504 -31678 377782 -24769 0 irq
rlabel metal1 s 369451 -13575 377901 -8217 0 VSS
rlabel metal1 s -117320 245880 -107876 253893 0 gpio<12>
rlabel metal1 s -117455 229677 -107460 236387 0 gpio<13>
rlabel metal1 s -117455 212877 -107460 219587 0 gpio<14>
rlabel metal1 s -117312 196029 -107603 203168 0 gpio<15>
rlabel metal1 s -117641 273192 -108233 279730 0 VSS
rlabel metal1 s -116217 290579 -108447 296323 0 VDD3V3
rlabel metal1 s -73117 315671 -66660 323257 0 gpio<10>
rlabel metal1 s -56317 315671 -49860 323257 0 gpio<9>
rlabel metal1 s -39517 315671 -33060 323257 0 gpio<8>
rlabel metal1 s -22717 315671 -16260 323257 0 gpio<7>
rlabel metal1 s -5917 315671 540 323257 0 gpio<6>
rlabel metal1 s 10883 315671 17340 323257 0 gpio<5>
rlabel metal1 s -89307 314732 -82676 323657 0 gpio<11>
rlabel metal1 s 369053 289951 377601 296125 0 spi_sdi
rlabel metal1 s 344449 316120 350390 323174 0 VDD3V3
rlabel metal1 s 145129 315690 151586 323276 0 gpio<0>
rlabel metal1 s 111529 315690 117986 323276 0 gpio<2>
rlabel metal1 s 128329 315690 134786 323276 0 gpio<1>
rlabel metal1 s 84729 315690 91186 323276 0 gpio<3>
rlabel metal1 s 67929 315690 74386 323276 0 gpio<4>
rlabel metal1 s 304823 316062 310764 323116 0 VDD3V3
rlabel metal1 s 321623 316062 327564 323116 0 VSS
rlabel metal1 s 285132 317000 287427 321592 0 VDD3V3
rlabel metal1 s 218762 317000 221057 321592 0 VDD1V8
rlabel metal1 370002 256958 377759 262815 0 spi_csb
rlabel metal1 s 369211 240020 378076 246035 0 spi_sck
rlabel metal1 s 369053 223557 378234 229256 0 spi_sdo
rlabel metal1 s 368979 149924 377408 155403 0 ser_tx
rlabel metal1 s 369816 167810 376581 172461 0 ser_rx
rlabel metal1 s 369940 274803 376306 279297 0 VSS
rlabel metal1 s 368961 122718 377921 129374 0 VDD1V8
rlabel metal1 s 369393 106440 376581 111514 0 VSS
rlabel metal1 s -20650 -69433 -14256 -60528 0 VDD3V3FC
rlabel metal1 s -87393 -69600 -81084 -60847 0 SDO
rlabel metal1 s -70290 -69844 -63641 -61138 0 SDI
rlabel metal1 -54460 -69686 -46703 -60979 0 CSB
rlabel metal1 -37838 -69686 -30715 -61613 0 SCK
rlabel metal1 s 4145 -67471 6518 -62988 0 VDD3V3
rlabel metal1 s 70472 -67471 72977 -62856 0 VDD1V8
<< end >>
