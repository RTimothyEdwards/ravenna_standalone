magic
tech EFXH018D
magscale 1 2
timestamp 1565723183
<< mimcap >>
rect -24745 32210 -20745 32240
rect -24745 28270 -24715 32210
rect -20775 28270 -20745 32210
rect -24745 28240 -20745 28270
rect -20215 32210 -16215 32240
rect -20215 28270 -20185 32210
rect -16245 28270 -16215 32210
rect -20215 28240 -16215 28270
rect -15685 32210 -11685 32240
rect -15685 28270 -15655 32210
rect -11715 28270 -11685 32210
rect -15685 28240 -11685 28270
rect -11155 32210 -7155 32240
rect -11155 28270 -11125 32210
rect -7185 28270 -7155 32210
rect -11155 28240 -7155 28270
rect -6625 32210 -2625 32240
rect -6625 28270 -6595 32210
rect -2655 28270 -2625 32210
rect -6625 28240 -2625 28270
rect -2095 32210 1905 32240
rect -2095 28270 -2065 32210
rect 1875 28270 1905 32210
rect -2095 28240 1905 28270
rect 2435 32210 6435 32240
rect 2435 28270 2465 32210
rect 6405 28270 6435 32210
rect 2435 28240 6435 28270
rect 6965 32210 10965 32240
rect 6965 28270 6995 32210
rect 10935 28270 10965 32210
rect 6965 28240 10965 28270
rect 11495 32210 15495 32240
rect 11495 28270 11525 32210
rect 15465 28270 15495 32210
rect 11495 28240 15495 28270
rect 16025 32210 20025 32240
rect 16025 28270 16055 32210
rect 19995 28270 20025 32210
rect 16025 28240 20025 28270
rect 20555 32210 24555 32240
rect 20555 28270 20585 32210
rect 24525 28270 24555 32210
rect 20555 28240 24555 28270
rect -24745 27890 -20745 27920
rect -24745 23950 -24715 27890
rect -20775 23950 -20745 27890
rect -24745 23920 -20745 23950
rect -20215 27890 -16215 27920
rect -20215 23950 -20185 27890
rect -16245 23950 -16215 27890
rect -20215 23920 -16215 23950
rect -15685 27890 -11685 27920
rect -15685 23950 -15655 27890
rect -11715 23950 -11685 27890
rect -15685 23920 -11685 23950
rect -11155 27890 -7155 27920
rect -11155 23950 -11125 27890
rect -7185 23950 -7155 27890
rect -11155 23920 -7155 23950
rect -6625 27890 -2625 27920
rect -6625 23950 -6595 27890
rect -2655 23950 -2625 27890
rect -6625 23920 -2625 23950
rect -2095 27890 1905 27920
rect -2095 23950 -2065 27890
rect 1875 23950 1905 27890
rect -2095 23920 1905 23950
rect 2435 27890 6435 27920
rect 2435 23950 2465 27890
rect 6405 23950 6435 27890
rect 2435 23920 6435 23950
rect 6965 27890 10965 27920
rect 6965 23950 6995 27890
rect 10935 23950 10965 27890
rect 6965 23920 10965 23950
rect 11495 27890 15495 27920
rect 11495 23950 11525 27890
rect 15465 23950 15495 27890
rect 11495 23920 15495 23950
rect 16025 27890 20025 27920
rect 16025 23950 16055 27890
rect 19995 23950 20025 27890
rect 16025 23920 20025 23950
rect 20555 27890 24555 27920
rect 20555 23950 20585 27890
rect 24525 23950 24555 27890
rect 20555 23920 24555 23950
rect -24745 23570 -20745 23600
rect -24745 19630 -24715 23570
rect -20775 19630 -20745 23570
rect -24745 19600 -20745 19630
rect -20215 23570 -16215 23600
rect -20215 19630 -20185 23570
rect -16245 19630 -16215 23570
rect -20215 19600 -16215 19630
rect -15685 23570 -11685 23600
rect -15685 19630 -15655 23570
rect -11715 19630 -11685 23570
rect -15685 19600 -11685 19630
rect -11155 23570 -7155 23600
rect -11155 19630 -11125 23570
rect -7185 19630 -7155 23570
rect -11155 19600 -7155 19630
rect -6625 23570 -2625 23600
rect -6625 19630 -6595 23570
rect -2655 19630 -2625 23570
rect -6625 19600 -2625 19630
rect -2095 23570 1905 23600
rect -2095 19630 -2065 23570
rect 1875 19630 1905 23570
rect -2095 19600 1905 19630
rect 2435 23570 6435 23600
rect 2435 19630 2465 23570
rect 6405 19630 6435 23570
rect 2435 19600 6435 19630
rect 6965 23570 10965 23600
rect 6965 19630 6995 23570
rect 10935 19630 10965 23570
rect 6965 19600 10965 19630
rect 11495 23570 15495 23600
rect 11495 19630 11525 23570
rect 15465 19630 15495 23570
rect 11495 19600 15495 19630
rect 16025 23570 20025 23600
rect 16025 19630 16055 23570
rect 19995 19630 20025 23570
rect 16025 19600 20025 19630
rect 20555 23570 24555 23600
rect 20555 19630 20585 23570
rect 24525 19630 24555 23570
rect 20555 19600 24555 19630
rect -24745 19250 -20745 19280
rect -24745 15310 -24715 19250
rect -20775 15310 -20745 19250
rect -24745 15280 -20745 15310
rect -20215 19250 -16215 19280
rect -20215 15310 -20185 19250
rect -16245 15310 -16215 19250
rect -20215 15280 -16215 15310
rect -15685 19250 -11685 19280
rect -15685 15310 -15655 19250
rect -11715 15310 -11685 19250
rect -15685 15280 -11685 15310
rect -11155 19250 -7155 19280
rect -11155 15310 -11125 19250
rect -7185 15310 -7155 19250
rect -11155 15280 -7155 15310
rect -6625 19250 -2625 19280
rect -6625 15310 -6595 19250
rect -2655 15310 -2625 19250
rect -6625 15280 -2625 15310
rect -2095 19250 1905 19280
rect -2095 15310 -2065 19250
rect 1875 15310 1905 19250
rect -2095 15280 1905 15310
rect 2435 19250 6435 19280
rect 2435 15310 2465 19250
rect 6405 15310 6435 19250
rect 2435 15280 6435 15310
rect 6965 19250 10965 19280
rect 6965 15310 6995 19250
rect 10935 15310 10965 19250
rect 6965 15280 10965 15310
rect 11495 19250 15495 19280
rect 11495 15310 11525 19250
rect 15465 15310 15495 19250
rect 11495 15280 15495 15310
rect 16025 19250 20025 19280
rect 16025 15310 16055 19250
rect 19995 15310 20025 19250
rect 16025 15280 20025 15310
rect 20555 19250 24555 19280
rect 20555 15310 20585 19250
rect 24525 15310 24555 19250
rect 20555 15280 24555 15310
rect -24745 14930 -20745 14960
rect -24745 10990 -24715 14930
rect -20775 10990 -20745 14930
rect -24745 10960 -20745 10990
rect -20215 14930 -16215 14960
rect -20215 10990 -20185 14930
rect -16245 10990 -16215 14930
rect -20215 10960 -16215 10990
rect -15685 14930 -11685 14960
rect -15685 10990 -15655 14930
rect -11715 10990 -11685 14930
rect -15685 10960 -11685 10990
rect -11155 14930 -7155 14960
rect -11155 10990 -11125 14930
rect -7185 10990 -7155 14930
rect -11155 10960 -7155 10990
rect -6625 14930 -2625 14960
rect -6625 10990 -6595 14930
rect -2655 10990 -2625 14930
rect -6625 10960 -2625 10990
rect -2095 14930 1905 14960
rect -2095 10990 -2065 14930
rect 1875 10990 1905 14930
rect -2095 10960 1905 10990
rect 2435 14930 6435 14960
rect 2435 10990 2465 14930
rect 6405 10990 6435 14930
rect 2435 10960 6435 10990
rect 6965 14930 10965 14960
rect 6965 10990 6995 14930
rect 10935 10990 10965 14930
rect 6965 10960 10965 10990
rect 11495 14930 15495 14960
rect 11495 10990 11525 14930
rect 15465 10990 15495 14930
rect 11495 10960 15495 10990
rect 16025 14930 20025 14960
rect 16025 10990 16055 14930
rect 19995 10990 20025 14930
rect 16025 10960 20025 10990
rect 20555 14930 24555 14960
rect 20555 10990 20585 14930
rect 24525 10990 24555 14930
rect 20555 10960 24555 10990
rect -24745 10610 -20745 10640
rect -24745 6670 -24715 10610
rect -20775 6670 -20745 10610
rect -24745 6640 -20745 6670
rect -20215 10610 -16215 10640
rect -20215 6670 -20185 10610
rect -16245 6670 -16215 10610
rect -20215 6640 -16215 6670
rect -15685 10610 -11685 10640
rect -15685 6670 -15655 10610
rect -11715 6670 -11685 10610
rect -15685 6640 -11685 6670
rect -11155 10610 -7155 10640
rect -11155 6670 -11125 10610
rect -7185 6670 -7155 10610
rect -11155 6640 -7155 6670
rect -6625 10610 -2625 10640
rect -6625 6670 -6595 10610
rect -2655 6670 -2625 10610
rect -6625 6640 -2625 6670
rect -2095 10610 1905 10640
rect -2095 6670 -2065 10610
rect 1875 6670 1905 10610
rect -2095 6640 1905 6670
rect 2435 10610 6435 10640
rect 2435 6670 2465 10610
rect 6405 6670 6435 10610
rect 2435 6640 6435 6670
rect 6965 10610 10965 10640
rect 6965 6670 6995 10610
rect 10935 6670 10965 10610
rect 6965 6640 10965 6670
rect 11495 10610 15495 10640
rect 11495 6670 11525 10610
rect 15465 6670 15495 10610
rect 11495 6640 15495 6670
rect 16025 10610 20025 10640
rect 16025 6670 16055 10610
rect 19995 6670 20025 10610
rect 16025 6640 20025 6670
rect 20555 10610 24555 10640
rect 20555 6670 20585 10610
rect 24525 6670 24555 10610
rect 20555 6640 24555 6670
rect -24745 6290 -20745 6320
rect -24745 2350 -24715 6290
rect -20775 2350 -20745 6290
rect -24745 2320 -20745 2350
rect -20215 6290 -16215 6320
rect -20215 2350 -20185 6290
rect -16245 2350 -16215 6290
rect -20215 2320 -16215 2350
rect -15685 6290 -11685 6320
rect -15685 2350 -15655 6290
rect -11715 2350 -11685 6290
rect -15685 2320 -11685 2350
rect -11155 6290 -7155 6320
rect -11155 2350 -11125 6290
rect -7185 2350 -7155 6290
rect -11155 2320 -7155 2350
rect -6625 6290 -2625 6320
rect -6625 2350 -6595 6290
rect -2655 2350 -2625 6290
rect -6625 2320 -2625 2350
rect -2095 6290 1905 6320
rect -2095 2350 -2065 6290
rect 1875 2350 1905 6290
rect -2095 2320 1905 2350
rect 2435 6290 6435 6320
rect 2435 2350 2465 6290
rect 6405 2350 6435 6290
rect 2435 2320 6435 2350
rect 6965 6290 10965 6320
rect 6965 2350 6995 6290
rect 10935 2350 10965 6290
rect 6965 2320 10965 2350
rect 11495 6290 15495 6320
rect 11495 2350 11525 6290
rect 15465 2350 15495 6290
rect 11495 2320 15495 2350
rect 16025 6290 20025 6320
rect 16025 2350 16055 6290
rect 19995 2350 20025 6290
rect 16025 2320 20025 2350
rect 20555 6290 24555 6320
rect 20555 2350 20585 6290
rect 24525 2350 24555 6290
rect 20555 2320 24555 2350
rect -24745 1970 -20745 2000
rect -24745 -1970 -24715 1970
rect -20775 -1970 -20745 1970
rect -24745 -2000 -20745 -1970
rect -20215 1970 -16215 2000
rect -20215 -1970 -20185 1970
rect -16245 -1970 -16215 1970
rect -20215 -2000 -16215 -1970
rect -15685 1970 -11685 2000
rect -15685 -1970 -15655 1970
rect -11715 -1970 -11685 1970
rect -15685 -2000 -11685 -1970
rect -11155 1970 -7155 2000
rect -11155 -1970 -11125 1970
rect -7185 -1970 -7155 1970
rect -11155 -2000 -7155 -1970
rect -6625 1970 -2625 2000
rect -6625 -1970 -6595 1970
rect -2655 -1970 -2625 1970
rect -6625 -2000 -2625 -1970
rect -2095 1970 1905 2000
rect -2095 -1970 -2065 1970
rect 1875 -1970 1905 1970
rect -2095 -2000 1905 -1970
rect 2435 1970 6435 2000
rect 2435 -1970 2465 1970
rect 6405 -1970 6435 1970
rect 2435 -2000 6435 -1970
rect 6965 1970 10965 2000
rect 6965 -1970 6995 1970
rect 10935 -1970 10965 1970
rect 6965 -2000 10965 -1970
rect 11495 1970 15495 2000
rect 11495 -1970 11525 1970
rect 15465 -1970 15495 1970
rect 11495 -2000 15495 -1970
rect 16025 1970 20025 2000
rect 16025 -1970 16055 1970
rect 19995 -1970 20025 1970
rect 16025 -2000 20025 -1970
rect 20555 1970 24555 2000
rect 20555 -1970 20585 1970
rect 24525 -1970 24555 1970
rect 20555 -2000 24555 -1970
rect -24745 -2350 -20745 -2320
rect -24745 -6290 -24715 -2350
rect -20775 -6290 -20745 -2350
rect -24745 -6320 -20745 -6290
rect -20215 -2350 -16215 -2320
rect -20215 -6290 -20185 -2350
rect -16245 -6290 -16215 -2350
rect -20215 -6320 -16215 -6290
rect -15685 -2350 -11685 -2320
rect -15685 -6290 -15655 -2350
rect -11715 -6290 -11685 -2350
rect -15685 -6320 -11685 -6290
rect -11155 -2350 -7155 -2320
rect -11155 -6290 -11125 -2350
rect -7185 -6290 -7155 -2350
rect -11155 -6320 -7155 -6290
rect -6625 -2350 -2625 -2320
rect -6625 -6290 -6595 -2350
rect -2655 -6290 -2625 -2350
rect -6625 -6320 -2625 -6290
rect -2095 -2350 1905 -2320
rect -2095 -6290 -2065 -2350
rect 1875 -6290 1905 -2350
rect -2095 -6320 1905 -6290
rect 2435 -2350 6435 -2320
rect 2435 -6290 2465 -2350
rect 6405 -6290 6435 -2350
rect 2435 -6320 6435 -6290
rect 6965 -2350 10965 -2320
rect 6965 -6290 6995 -2350
rect 10935 -6290 10965 -2350
rect 6965 -6320 10965 -6290
rect 11495 -2350 15495 -2320
rect 11495 -6290 11525 -2350
rect 15465 -6290 15495 -2350
rect 11495 -6320 15495 -6290
rect 16025 -2350 20025 -2320
rect 16025 -6290 16055 -2350
rect 19995 -6290 20025 -2350
rect 16025 -6320 20025 -6290
rect 20555 -2350 24555 -2320
rect 20555 -6290 20585 -2350
rect 24525 -6290 24555 -2350
rect 20555 -6320 24555 -6290
rect -24745 -6670 -20745 -6640
rect -24745 -10610 -24715 -6670
rect -20775 -10610 -20745 -6670
rect -24745 -10640 -20745 -10610
rect -20215 -6670 -16215 -6640
rect -20215 -10610 -20185 -6670
rect -16245 -10610 -16215 -6670
rect -20215 -10640 -16215 -10610
rect -15685 -6670 -11685 -6640
rect -15685 -10610 -15655 -6670
rect -11715 -10610 -11685 -6670
rect -15685 -10640 -11685 -10610
rect -11155 -6670 -7155 -6640
rect -11155 -10610 -11125 -6670
rect -7185 -10610 -7155 -6670
rect -11155 -10640 -7155 -10610
rect -6625 -6670 -2625 -6640
rect -6625 -10610 -6595 -6670
rect -2655 -10610 -2625 -6670
rect -6625 -10640 -2625 -10610
rect -2095 -6670 1905 -6640
rect -2095 -10610 -2065 -6670
rect 1875 -10610 1905 -6670
rect -2095 -10640 1905 -10610
rect 2435 -6670 6435 -6640
rect 2435 -10610 2465 -6670
rect 6405 -10610 6435 -6670
rect 2435 -10640 6435 -10610
rect 6965 -6670 10965 -6640
rect 6965 -10610 6995 -6670
rect 10935 -10610 10965 -6670
rect 6965 -10640 10965 -10610
rect 11495 -6670 15495 -6640
rect 11495 -10610 11525 -6670
rect 15465 -10610 15495 -6670
rect 11495 -10640 15495 -10610
rect 16025 -6670 20025 -6640
rect 16025 -10610 16055 -6670
rect 19995 -10610 20025 -6670
rect 16025 -10640 20025 -10610
rect 20555 -6670 24555 -6640
rect 20555 -10610 20585 -6670
rect 24525 -10610 24555 -6670
rect 20555 -10640 24555 -10610
rect -24745 -10990 -20745 -10960
rect -24745 -14930 -24715 -10990
rect -20775 -14930 -20745 -10990
rect -24745 -14960 -20745 -14930
rect -20215 -10990 -16215 -10960
rect -20215 -14930 -20185 -10990
rect -16245 -14930 -16215 -10990
rect -20215 -14960 -16215 -14930
rect -15685 -10990 -11685 -10960
rect -15685 -14930 -15655 -10990
rect -11715 -14930 -11685 -10990
rect -15685 -14960 -11685 -14930
rect -11155 -10990 -7155 -10960
rect -11155 -14930 -11125 -10990
rect -7185 -14930 -7155 -10990
rect -11155 -14960 -7155 -14930
rect -6625 -10990 -2625 -10960
rect -6625 -14930 -6595 -10990
rect -2655 -14930 -2625 -10990
rect -6625 -14960 -2625 -14930
rect -2095 -10990 1905 -10960
rect -2095 -14930 -2065 -10990
rect 1875 -14930 1905 -10990
rect -2095 -14960 1905 -14930
rect 2435 -10990 6435 -10960
rect 2435 -14930 2465 -10990
rect 6405 -14930 6435 -10990
rect 2435 -14960 6435 -14930
rect 6965 -10990 10965 -10960
rect 6965 -14930 6995 -10990
rect 10935 -14930 10965 -10990
rect 6965 -14960 10965 -14930
rect 11495 -10990 15495 -10960
rect 11495 -14930 11525 -10990
rect 15465 -14930 15495 -10990
rect 11495 -14960 15495 -14930
rect 16025 -10990 20025 -10960
rect 16025 -14930 16055 -10990
rect 19995 -14930 20025 -10990
rect 16025 -14960 20025 -14930
rect 20555 -10990 24555 -10960
rect 20555 -14930 20585 -10990
rect 24525 -14930 24555 -10990
rect 20555 -14960 24555 -14930
rect -24745 -15310 -20745 -15280
rect -24745 -19250 -24715 -15310
rect -20775 -19250 -20745 -15310
rect -24745 -19280 -20745 -19250
rect -20215 -15310 -16215 -15280
rect -20215 -19250 -20185 -15310
rect -16245 -19250 -16215 -15310
rect -20215 -19280 -16215 -19250
rect -15685 -15310 -11685 -15280
rect -15685 -19250 -15655 -15310
rect -11715 -19250 -11685 -15310
rect -15685 -19280 -11685 -19250
rect -11155 -15310 -7155 -15280
rect -11155 -19250 -11125 -15310
rect -7185 -19250 -7155 -15310
rect -11155 -19280 -7155 -19250
rect -6625 -15310 -2625 -15280
rect -6625 -19250 -6595 -15310
rect -2655 -19250 -2625 -15310
rect -6625 -19280 -2625 -19250
rect -2095 -15310 1905 -15280
rect -2095 -19250 -2065 -15310
rect 1875 -19250 1905 -15310
rect -2095 -19280 1905 -19250
rect 2435 -15310 6435 -15280
rect 2435 -19250 2465 -15310
rect 6405 -19250 6435 -15310
rect 2435 -19280 6435 -19250
rect 6965 -15310 10965 -15280
rect 6965 -19250 6995 -15310
rect 10935 -19250 10965 -15310
rect 6965 -19280 10965 -19250
rect 11495 -15310 15495 -15280
rect 11495 -19250 11525 -15310
rect 15465 -19250 15495 -15310
rect 11495 -19280 15495 -19250
rect 16025 -15310 20025 -15280
rect 16025 -19250 16055 -15310
rect 19995 -19250 20025 -15310
rect 16025 -19280 20025 -19250
rect 20555 -15310 24555 -15280
rect 20555 -19250 20585 -15310
rect 24525 -19250 24555 -15310
rect 20555 -19280 24555 -19250
rect -24745 -19630 -20745 -19600
rect -24745 -23570 -24715 -19630
rect -20775 -23570 -20745 -19630
rect -24745 -23600 -20745 -23570
rect -20215 -19630 -16215 -19600
rect -20215 -23570 -20185 -19630
rect -16245 -23570 -16215 -19630
rect -20215 -23600 -16215 -23570
rect -15685 -19630 -11685 -19600
rect -15685 -23570 -15655 -19630
rect -11715 -23570 -11685 -19630
rect -15685 -23600 -11685 -23570
rect -11155 -19630 -7155 -19600
rect -11155 -23570 -11125 -19630
rect -7185 -23570 -7155 -19630
rect -11155 -23600 -7155 -23570
rect -6625 -19630 -2625 -19600
rect -6625 -23570 -6595 -19630
rect -2655 -23570 -2625 -19630
rect -6625 -23600 -2625 -23570
rect -2095 -19630 1905 -19600
rect -2095 -23570 -2065 -19630
rect 1875 -23570 1905 -19630
rect -2095 -23600 1905 -23570
rect 2435 -19630 6435 -19600
rect 2435 -23570 2465 -19630
rect 6405 -23570 6435 -19630
rect 2435 -23600 6435 -23570
rect 6965 -19630 10965 -19600
rect 6965 -23570 6995 -19630
rect 10935 -23570 10965 -19630
rect 6965 -23600 10965 -23570
rect 11495 -19630 15495 -19600
rect 11495 -23570 11525 -19630
rect 15465 -23570 15495 -19630
rect 11495 -23600 15495 -23570
rect 16025 -19630 20025 -19600
rect 16025 -23570 16055 -19630
rect 19995 -23570 20025 -19630
rect 16025 -23600 20025 -23570
rect 20555 -19630 24555 -19600
rect 20555 -23570 20585 -19630
rect 24525 -23570 24555 -19630
rect 20555 -23600 24555 -23570
rect -24745 -23950 -20745 -23920
rect -24745 -27890 -24715 -23950
rect -20775 -27890 -20745 -23950
rect -24745 -27920 -20745 -27890
rect -20215 -23950 -16215 -23920
rect -20215 -27890 -20185 -23950
rect -16245 -27890 -16215 -23950
rect -20215 -27920 -16215 -27890
rect -15685 -23950 -11685 -23920
rect -15685 -27890 -15655 -23950
rect -11715 -27890 -11685 -23950
rect -15685 -27920 -11685 -27890
rect -11155 -23950 -7155 -23920
rect -11155 -27890 -11125 -23950
rect -7185 -27890 -7155 -23950
rect -11155 -27920 -7155 -27890
rect -6625 -23950 -2625 -23920
rect -6625 -27890 -6595 -23950
rect -2655 -27890 -2625 -23950
rect -6625 -27920 -2625 -27890
rect -2095 -23950 1905 -23920
rect -2095 -27890 -2065 -23950
rect 1875 -27890 1905 -23950
rect -2095 -27920 1905 -27890
rect 2435 -23950 6435 -23920
rect 2435 -27890 2465 -23950
rect 6405 -27890 6435 -23950
rect 2435 -27920 6435 -27890
rect 6965 -23950 10965 -23920
rect 6965 -27890 6995 -23950
rect 10935 -27890 10965 -23950
rect 6965 -27920 10965 -27890
rect 11495 -23950 15495 -23920
rect 11495 -27890 11525 -23950
rect 15465 -27890 15495 -23950
rect 11495 -27920 15495 -27890
rect 16025 -23950 20025 -23920
rect 16025 -27890 16055 -23950
rect 19995 -27890 20025 -23950
rect 16025 -27920 20025 -27890
rect 20555 -23950 24555 -23920
rect 20555 -27890 20585 -23950
rect 24525 -27890 24555 -23950
rect 20555 -27920 24555 -27890
rect -24745 -28270 -20745 -28240
rect -24745 -32210 -24715 -28270
rect -20775 -32210 -20745 -28270
rect -24745 -32240 -20745 -32210
rect -20215 -28270 -16215 -28240
rect -20215 -32210 -20185 -28270
rect -16245 -32210 -16215 -28270
rect -20215 -32240 -16215 -32210
rect -15685 -28270 -11685 -28240
rect -15685 -32210 -15655 -28270
rect -11715 -32210 -11685 -28270
rect -15685 -32240 -11685 -32210
rect -11155 -28270 -7155 -28240
rect -11155 -32210 -11125 -28270
rect -7185 -32210 -7155 -28270
rect -11155 -32240 -7155 -32210
rect -6625 -28270 -2625 -28240
rect -6625 -32210 -6595 -28270
rect -2655 -32210 -2625 -28270
rect -6625 -32240 -2625 -32210
rect -2095 -28270 1905 -28240
rect -2095 -32210 -2065 -28270
rect 1875 -32210 1905 -28270
rect -2095 -32240 1905 -32210
rect 2435 -28270 6435 -28240
rect 2435 -32210 2465 -28270
rect 6405 -32210 6435 -28270
rect 2435 -32240 6435 -32210
rect 6965 -28270 10965 -28240
rect 6965 -32210 6995 -28270
rect 10935 -32210 10965 -28270
rect 6965 -32240 10965 -32210
rect 11495 -28270 15495 -28240
rect 11495 -32210 11525 -28270
rect 15465 -32210 15495 -28270
rect 11495 -32240 15495 -32210
rect 16025 -28270 20025 -28240
rect 16025 -32210 16055 -28270
rect 19995 -32210 20025 -28270
rect 16025 -32240 20025 -32210
rect 20555 -28270 24555 -28240
rect 20555 -32210 20585 -28270
rect 24525 -32210 24555 -28270
rect 20555 -32240 24555 -32210
<< mimcapcontact >>
rect -24715 28270 -20775 32210
rect -20185 28270 -16245 32210
rect -15655 28270 -11715 32210
rect -11125 28270 -7185 32210
rect -6595 28270 -2655 32210
rect -2065 28270 1875 32210
rect 2465 28270 6405 32210
rect 6995 28270 10935 32210
rect 11525 28270 15465 32210
rect 16055 28270 19995 32210
rect 20585 28270 24525 32210
rect -24715 23950 -20775 27890
rect -20185 23950 -16245 27890
rect -15655 23950 -11715 27890
rect -11125 23950 -7185 27890
rect -6595 23950 -2655 27890
rect -2065 23950 1875 27890
rect 2465 23950 6405 27890
rect 6995 23950 10935 27890
rect 11525 23950 15465 27890
rect 16055 23950 19995 27890
rect 20585 23950 24525 27890
rect -24715 19630 -20775 23570
rect -20185 19630 -16245 23570
rect -15655 19630 -11715 23570
rect -11125 19630 -7185 23570
rect -6595 19630 -2655 23570
rect -2065 19630 1875 23570
rect 2465 19630 6405 23570
rect 6995 19630 10935 23570
rect 11525 19630 15465 23570
rect 16055 19630 19995 23570
rect 20585 19630 24525 23570
rect -24715 15310 -20775 19250
rect -20185 15310 -16245 19250
rect -15655 15310 -11715 19250
rect -11125 15310 -7185 19250
rect -6595 15310 -2655 19250
rect -2065 15310 1875 19250
rect 2465 15310 6405 19250
rect 6995 15310 10935 19250
rect 11525 15310 15465 19250
rect 16055 15310 19995 19250
rect 20585 15310 24525 19250
rect -24715 10990 -20775 14930
rect -20185 10990 -16245 14930
rect -15655 10990 -11715 14930
rect -11125 10990 -7185 14930
rect -6595 10990 -2655 14930
rect -2065 10990 1875 14930
rect 2465 10990 6405 14930
rect 6995 10990 10935 14930
rect 11525 10990 15465 14930
rect 16055 10990 19995 14930
rect 20585 10990 24525 14930
rect -24715 6670 -20775 10610
rect -20185 6670 -16245 10610
rect -15655 6670 -11715 10610
rect -11125 6670 -7185 10610
rect -6595 6670 -2655 10610
rect -2065 6670 1875 10610
rect 2465 6670 6405 10610
rect 6995 6670 10935 10610
rect 11525 6670 15465 10610
rect 16055 6670 19995 10610
rect 20585 6670 24525 10610
rect -24715 2350 -20775 6290
rect -20185 2350 -16245 6290
rect -15655 2350 -11715 6290
rect -11125 2350 -7185 6290
rect -6595 2350 -2655 6290
rect -2065 2350 1875 6290
rect 2465 2350 6405 6290
rect 6995 2350 10935 6290
rect 11525 2350 15465 6290
rect 16055 2350 19995 6290
rect 20585 2350 24525 6290
rect -24715 -1970 -20775 1970
rect -20185 -1970 -16245 1970
rect -15655 -1970 -11715 1970
rect -11125 -1970 -7185 1970
rect -6595 -1970 -2655 1970
rect -2065 -1970 1875 1970
rect 2465 -1970 6405 1970
rect 6995 -1970 10935 1970
rect 11525 -1970 15465 1970
rect 16055 -1970 19995 1970
rect 20585 -1970 24525 1970
rect -24715 -6290 -20775 -2350
rect -20185 -6290 -16245 -2350
rect -15655 -6290 -11715 -2350
rect -11125 -6290 -7185 -2350
rect -6595 -6290 -2655 -2350
rect -2065 -6290 1875 -2350
rect 2465 -6290 6405 -2350
rect 6995 -6290 10935 -2350
rect 11525 -6290 15465 -2350
rect 16055 -6290 19995 -2350
rect 20585 -6290 24525 -2350
rect -24715 -10610 -20775 -6670
rect -20185 -10610 -16245 -6670
rect -15655 -10610 -11715 -6670
rect -11125 -10610 -7185 -6670
rect -6595 -10610 -2655 -6670
rect -2065 -10610 1875 -6670
rect 2465 -10610 6405 -6670
rect 6995 -10610 10935 -6670
rect 11525 -10610 15465 -6670
rect 16055 -10610 19995 -6670
rect 20585 -10610 24525 -6670
rect -24715 -14930 -20775 -10990
rect -20185 -14930 -16245 -10990
rect -15655 -14930 -11715 -10990
rect -11125 -14930 -7185 -10990
rect -6595 -14930 -2655 -10990
rect -2065 -14930 1875 -10990
rect 2465 -14930 6405 -10990
rect 6995 -14930 10935 -10990
rect 11525 -14930 15465 -10990
rect 16055 -14930 19995 -10990
rect 20585 -14930 24525 -10990
rect -24715 -19250 -20775 -15310
rect -20185 -19250 -16245 -15310
rect -15655 -19250 -11715 -15310
rect -11125 -19250 -7185 -15310
rect -6595 -19250 -2655 -15310
rect -2065 -19250 1875 -15310
rect 2465 -19250 6405 -15310
rect 6995 -19250 10935 -15310
rect 11525 -19250 15465 -15310
rect 16055 -19250 19995 -15310
rect 20585 -19250 24525 -15310
rect -24715 -23570 -20775 -19630
rect -20185 -23570 -16245 -19630
rect -15655 -23570 -11715 -19630
rect -11125 -23570 -7185 -19630
rect -6595 -23570 -2655 -19630
rect -2065 -23570 1875 -19630
rect 2465 -23570 6405 -19630
rect 6995 -23570 10935 -19630
rect 11525 -23570 15465 -19630
rect 16055 -23570 19995 -19630
rect 20585 -23570 24525 -19630
rect -24715 -27890 -20775 -23950
rect -20185 -27890 -16245 -23950
rect -15655 -27890 -11715 -23950
rect -11125 -27890 -7185 -23950
rect -6595 -27890 -2655 -23950
rect -2065 -27890 1875 -23950
rect 2465 -27890 6405 -23950
rect 6995 -27890 10935 -23950
rect 11525 -27890 15465 -23950
rect 16055 -27890 19995 -23950
rect 20585 -27890 24525 -23950
rect -24715 -32210 -20775 -28270
rect -20185 -32210 -16245 -28270
rect -15655 -32210 -11715 -28270
rect -11125 -32210 -7185 -28270
rect -6595 -32210 -2655 -28270
rect -2065 -32210 1875 -28270
rect 2465 -32210 6405 -28270
rect 6995 -32210 10935 -28270
rect 11525 -32210 15465 -28270
rect 16055 -32210 19995 -28270
rect 20585 -32210 24525 -28270
<< metal4 >>
rect -24845 32312 -20455 32340
rect -24845 32240 -20575 32312
rect -24845 28240 -24745 32240
rect -20745 28240 -20575 32240
rect -24845 28168 -20575 28240
rect -20475 28168 -20455 32312
rect -24845 28140 -20455 28168
rect -20315 32312 -15925 32340
rect -20315 32240 -16045 32312
rect -20315 28240 -20215 32240
rect -16215 28240 -16045 32240
rect -20315 28168 -16045 28240
rect -15945 28168 -15925 32312
rect -20315 28140 -15925 28168
rect -15785 32312 -11395 32340
rect -15785 32240 -11515 32312
rect -15785 28240 -15685 32240
rect -11685 28240 -11515 32240
rect -15785 28168 -11515 28240
rect -11415 28168 -11395 32312
rect -15785 28140 -11395 28168
rect -11255 32312 -6865 32340
rect -11255 32240 -6985 32312
rect -11255 28240 -11155 32240
rect -7155 28240 -6985 32240
rect -11255 28168 -6985 28240
rect -6885 28168 -6865 32312
rect -11255 28140 -6865 28168
rect -6725 32312 -2335 32340
rect -6725 32240 -2455 32312
rect -6725 28240 -6625 32240
rect -2625 28240 -2455 32240
rect -6725 28168 -2455 28240
rect -2355 28168 -2335 32312
rect -6725 28140 -2335 28168
rect -2195 32312 2195 32340
rect -2195 32240 2075 32312
rect -2195 28240 -2095 32240
rect 1905 28240 2075 32240
rect -2195 28168 2075 28240
rect 2175 28168 2195 32312
rect -2195 28140 2195 28168
rect 2335 32312 6725 32340
rect 2335 32240 6605 32312
rect 2335 28240 2435 32240
rect 6435 28240 6605 32240
rect 2335 28168 6605 28240
rect 6705 28168 6725 32312
rect 2335 28140 6725 28168
rect 6865 32312 11255 32340
rect 6865 32240 11135 32312
rect 6865 28240 6965 32240
rect 10965 28240 11135 32240
rect 6865 28168 11135 28240
rect 11235 28168 11255 32312
rect 6865 28140 11255 28168
rect 11395 32312 15785 32340
rect 11395 32240 15665 32312
rect 11395 28240 11495 32240
rect 15495 28240 15665 32240
rect 11395 28168 15665 28240
rect 15765 28168 15785 32312
rect 11395 28140 15785 28168
rect 15925 32312 20315 32340
rect 15925 32240 20195 32312
rect 15925 28240 16025 32240
rect 20025 28240 20195 32240
rect 15925 28168 20195 28240
rect 20295 28168 20315 32312
rect 15925 28140 20315 28168
rect 20455 32312 24845 32340
rect 20455 32240 24725 32312
rect 20455 28240 20555 32240
rect 24555 28240 24725 32240
rect 20455 28168 24725 28240
rect 24825 28168 24845 32312
rect 20455 28140 24845 28168
rect -24845 27992 -20455 28020
rect -24845 27920 -20575 27992
rect -24845 23920 -24745 27920
rect -20745 23920 -20575 27920
rect -24845 23848 -20575 23920
rect -20475 23848 -20455 27992
rect -24845 23820 -20455 23848
rect -20315 27992 -15925 28020
rect -20315 27920 -16045 27992
rect -20315 23920 -20215 27920
rect -16215 23920 -16045 27920
rect -20315 23848 -16045 23920
rect -15945 23848 -15925 27992
rect -20315 23820 -15925 23848
rect -15785 27992 -11395 28020
rect -15785 27920 -11515 27992
rect -15785 23920 -15685 27920
rect -11685 23920 -11515 27920
rect -15785 23848 -11515 23920
rect -11415 23848 -11395 27992
rect -15785 23820 -11395 23848
rect -11255 27992 -6865 28020
rect -11255 27920 -6985 27992
rect -11255 23920 -11155 27920
rect -7155 23920 -6985 27920
rect -11255 23848 -6985 23920
rect -6885 23848 -6865 27992
rect -11255 23820 -6865 23848
rect -6725 27992 -2335 28020
rect -6725 27920 -2455 27992
rect -6725 23920 -6625 27920
rect -2625 23920 -2455 27920
rect -6725 23848 -2455 23920
rect -2355 23848 -2335 27992
rect -6725 23820 -2335 23848
rect -2195 27992 2195 28020
rect -2195 27920 2075 27992
rect -2195 23920 -2095 27920
rect 1905 23920 2075 27920
rect -2195 23848 2075 23920
rect 2175 23848 2195 27992
rect -2195 23820 2195 23848
rect 2335 27992 6725 28020
rect 2335 27920 6605 27992
rect 2335 23920 2435 27920
rect 6435 23920 6605 27920
rect 2335 23848 6605 23920
rect 6705 23848 6725 27992
rect 2335 23820 6725 23848
rect 6865 27992 11255 28020
rect 6865 27920 11135 27992
rect 6865 23920 6965 27920
rect 10965 23920 11135 27920
rect 6865 23848 11135 23920
rect 11235 23848 11255 27992
rect 6865 23820 11255 23848
rect 11395 27992 15785 28020
rect 11395 27920 15665 27992
rect 11395 23920 11495 27920
rect 15495 23920 15665 27920
rect 11395 23848 15665 23920
rect 15765 23848 15785 27992
rect 11395 23820 15785 23848
rect 15925 27992 20315 28020
rect 15925 27920 20195 27992
rect 15925 23920 16025 27920
rect 20025 23920 20195 27920
rect 15925 23848 20195 23920
rect 20295 23848 20315 27992
rect 15925 23820 20315 23848
rect 20455 27992 24845 28020
rect 20455 27920 24725 27992
rect 20455 23920 20555 27920
rect 24555 23920 24725 27920
rect 20455 23848 24725 23920
rect 24825 23848 24845 27992
rect 20455 23820 24845 23848
rect -24845 23672 -20455 23700
rect -24845 23600 -20575 23672
rect -24845 19600 -24745 23600
rect -20745 19600 -20575 23600
rect -24845 19528 -20575 19600
rect -20475 19528 -20455 23672
rect -24845 19500 -20455 19528
rect -20315 23672 -15925 23700
rect -20315 23600 -16045 23672
rect -20315 19600 -20215 23600
rect -16215 19600 -16045 23600
rect -20315 19528 -16045 19600
rect -15945 19528 -15925 23672
rect -20315 19500 -15925 19528
rect -15785 23672 -11395 23700
rect -15785 23600 -11515 23672
rect -15785 19600 -15685 23600
rect -11685 19600 -11515 23600
rect -15785 19528 -11515 19600
rect -11415 19528 -11395 23672
rect -15785 19500 -11395 19528
rect -11255 23672 -6865 23700
rect -11255 23600 -6985 23672
rect -11255 19600 -11155 23600
rect -7155 19600 -6985 23600
rect -11255 19528 -6985 19600
rect -6885 19528 -6865 23672
rect -11255 19500 -6865 19528
rect -6725 23672 -2335 23700
rect -6725 23600 -2455 23672
rect -6725 19600 -6625 23600
rect -2625 19600 -2455 23600
rect -6725 19528 -2455 19600
rect -2355 19528 -2335 23672
rect -6725 19500 -2335 19528
rect -2195 23672 2195 23700
rect -2195 23600 2075 23672
rect -2195 19600 -2095 23600
rect 1905 19600 2075 23600
rect -2195 19528 2075 19600
rect 2175 19528 2195 23672
rect -2195 19500 2195 19528
rect 2335 23672 6725 23700
rect 2335 23600 6605 23672
rect 2335 19600 2435 23600
rect 6435 19600 6605 23600
rect 2335 19528 6605 19600
rect 6705 19528 6725 23672
rect 2335 19500 6725 19528
rect 6865 23672 11255 23700
rect 6865 23600 11135 23672
rect 6865 19600 6965 23600
rect 10965 19600 11135 23600
rect 6865 19528 11135 19600
rect 11235 19528 11255 23672
rect 6865 19500 11255 19528
rect 11395 23672 15785 23700
rect 11395 23600 15665 23672
rect 11395 19600 11495 23600
rect 15495 19600 15665 23600
rect 11395 19528 15665 19600
rect 15765 19528 15785 23672
rect 11395 19500 15785 19528
rect 15925 23672 20315 23700
rect 15925 23600 20195 23672
rect 15925 19600 16025 23600
rect 20025 19600 20195 23600
rect 15925 19528 20195 19600
rect 20295 19528 20315 23672
rect 15925 19500 20315 19528
rect 20455 23672 24845 23700
rect 20455 23600 24725 23672
rect 20455 19600 20555 23600
rect 24555 19600 24725 23600
rect 20455 19528 24725 19600
rect 24825 19528 24845 23672
rect 20455 19500 24845 19528
rect -24845 19352 -20455 19380
rect -24845 19280 -20575 19352
rect -24845 15280 -24745 19280
rect -20745 15280 -20575 19280
rect -24845 15208 -20575 15280
rect -20475 15208 -20455 19352
rect -24845 15180 -20455 15208
rect -20315 19352 -15925 19380
rect -20315 19280 -16045 19352
rect -20315 15280 -20215 19280
rect -16215 15280 -16045 19280
rect -20315 15208 -16045 15280
rect -15945 15208 -15925 19352
rect -20315 15180 -15925 15208
rect -15785 19352 -11395 19380
rect -15785 19280 -11515 19352
rect -15785 15280 -15685 19280
rect -11685 15280 -11515 19280
rect -15785 15208 -11515 15280
rect -11415 15208 -11395 19352
rect -15785 15180 -11395 15208
rect -11255 19352 -6865 19380
rect -11255 19280 -6985 19352
rect -11255 15280 -11155 19280
rect -7155 15280 -6985 19280
rect -11255 15208 -6985 15280
rect -6885 15208 -6865 19352
rect -11255 15180 -6865 15208
rect -6725 19352 -2335 19380
rect -6725 19280 -2455 19352
rect -6725 15280 -6625 19280
rect -2625 15280 -2455 19280
rect -6725 15208 -2455 15280
rect -2355 15208 -2335 19352
rect -6725 15180 -2335 15208
rect -2195 19352 2195 19380
rect -2195 19280 2075 19352
rect -2195 15280 -2095 19280
rect 1905 15280 2075 19280
rect -2195 15208 2075 15280
rect 2175 15208 2195 19352
rect -2195 15180 2195 15208
rect 2335 19352 6725 19380
rect 2335 19280 6605 19352
rect 2335 15280 2435 19280
rect 6435 15280 6605 19280
rect 2335 15208 6605 15280
rect 6705 15208 6725 19352
rect 2335 15180 6725 15208
rect 6865 19352 11255 19380
rect 6865 19280 11135 19352
rect 6865 15280 6965 19280
rect 10965 15280 11135 19280
rect 6865 15208 11135 15280
rect 11235 15208 11255 19352
rect 6865 15180 11255 15208
rect 11395 19352 15785 19380
rect 11395 19280 15665 19352
rect 11395 15280 11495 19280
rect 15495 15280 15665 19280
rect 11395 15208 15665 15280
rect 15765 15208 15785 19352
rect 11395 15180 15785 15208
rect 15925 19352 20315 19380
rect 15925 19280 20195 19352
rect 15925 15280 16025 19280
rect 20025 15280 20195 19280
rect 15925 15208 20195 15280
rect 20295 15208 20315 19352
rect 15925 15180 20315 15208
rect 20455 19352 24845 19380
rect 20455 19280 24725 19352
rect 20455 15280 20555 19280
rect 24555 15280 24725 19280
rect 20455 15208 24725 15280
rect 24825 15208 24845 19352
rect 20455 15180 24845 15208
rect -24845 15032 -20455 15060
rect -24845 14960 -20575 15032
rect -24845 10960 -24745 14960
rect -20745 10960 -20575 14960
rect -24845 10888 -20575 10960
rect -20475 10888 -20455 15032
rect -24845 10860 -20455 10888
rect -20315 15032 -15925 15060
rect -20315 14960 -16045 15032
rect -20315 10960 -20215 14960
rect -16215 10960 -16045 14960
rect -20315 10888 -16045 10960
rect -15945 10888 -15925 15032
rect -20315 10860 -15925 10888
rect -15785 15032 -11395 15060
rect -15785 14960 -11515 15032
rect -15785 10960 -15685 14960
rect -11685 10960 -11515 14960
rect -15785 10888 -11515 10960
rect -11415 10888 -11395 15032
rect -15785 10860 -11395 10888
rect -11255 15032 -6865 15060
rect -11255 14960 -6985 15032
rect -11255 10960 -11155 14960
rect -7155 10960 -6985 14960
rect -11255 10888 -6985 10960
rect -6885 10888 -6865 15032
rect -11255 10860 -6865 10888
rect -6725 15032 -2335 15060
rect -6725 14960 -2455 15032
rect -6725 10960 -6625 14960
rect -2625 10960 -2455 14960
rect -6725 10888 -2455 10960
rect -2355 10888 -2335 15032
rect -6725 10860 -2335 10888
rect -2195 15032 2195 15060
rect -2195 14960 2075 15032
rect -2195 10960 -2095 14960
rect 1905 10960 2075 14960
rect -2195 10888 2075 10960
rect 2175 10888 2195 15032
rect -2195 10860 2195 10888
rect 2335 15032 6725 15060
rect 2335 14960 6605 15032
rect 2335 10960 2435 14960
rect 6435 10960 6605 14960
rect 2335 10888 6605 10960
rect 6705 10888 6725 15032
rect 2335 10860 6725 10888
rect 6865 15032 11255 15060
rect 6865 14960 11135 15032
rect 6865 10960 6965 14960
rect 10965 10960 11135 14960
rect 6865 10888 11135 10960
rect 11235 10888 11255 15032
rect 6865 10860 11255 10888
rect 11395 15032 15785 15060
rect 11395 14960 15665 15032
rect 11395 10960 11495 14960
rect 15495 10960 15665 14960
rect 11395 10888 15665 10960
rect 15765 10888 15785 15032
rect 11395 10860 15785 10888
rect 15925 15032 20315 15060
rect 15925 14960 20195 15032
rect 15925 10960 16025 14960
rect 20025 10960 20195 14960
rect 15925 10888 20195 10960
rect 20295 10888 20315 15032
rect 15925 10860 20315 10888
rect 20455 15032 24845 15060
rect 20455 14960 24725 15032
rect 20455 10960 20555 14960
rect 24555 10960 24725 14960
rect 20455 10888 24725 10960
rect 24825 10888 24845 15032
rect 20455 10860 24845 10888
rect -24845 10712 -20455 10740
rect -24845 10640 -20575 10712
rect -24845 6640 -24745 10640
rect -20745 6640 -20575 10640
rect -24845 6568 -20575 6640
rect -20475 6568 -20455 10712
rect -24845 6540 -20455 6568
rect -20315 10712 -15925 10740
rect -20315 10640 -16045 10712
rect -20315 6640 -20215 10640
rect -16215 6640 -16045 10640
rect -20315 6568 -16045 6640
rect -15945 6568 -15925 10712
rect -20315 6540 -15925 6568
rect -15785 10712 -11395 10740
rect -15785 10640 -11515 10712
rect -15785 6640 -15685 10640
rect -11685 6640 -11515 10640
rect -15785 6568 -11515 6640
rect -11415 6568 -11395 10712
rect -15785 6540 -11395 6568
rect -11255 10712 -6865 10740
rect -11255 10640 -6985 10712
rect -11255 6640 -11155 10640
rect -7155 6640 -6985 10640
rect -11255 6568 -6985 6640
rect -6885 6568 -6865 10712
rect -11255 6540 -6865 6568
rect -6725 10712 -2335 10740
rect -6725 10640 -2455 10712
rect -6725 6640 -6625 10640
rect -2625 6640 -2455 10640
rect -6725 6568 -2455 6640
rect -2355 6568 -2335 10712
rect -6725 6540 -2335 6568
rect -2195 10712 2195 10740
rect -2195 10640 2075 10712
rect -2195 6640 -2095 10640
rect 1905 6640 2075 10640
rect -2195 6568 2075 6640
rect 2175 6568 2195 10712
rect -2195 6540 2195 6568
rect 2335 10712 6725 10740
rect 2335 10640 6605 10712
rect 2335 6640 2435 10640
rect 6435 6640 6605 10640
rect 2335 6568 6605 6640
rect 6705 6568 6725 10712
rect 2335 6540 6725 6568
rect 6865 10712 11255 10740
rect 6865 10640 11135 10712
rect 6865 6640 6965 10640
rect 10965 6640 11135 10640
rect 6865 6568 11135 6640
rect 11235 6568 11255 10712
rect 6865 6540 11255 6568
rect 11395 10712 15785 10740
rect 11395 10640 15665 10712
rect 11395 6640 11495 10640
rect 15495 6640 15665 10640
rect 11395 6568 15665 6640
rect 15765 6568 15785 10712
rect 11395 6540 15785 6568
rect 15925 10712 20315 10740
rect 15925 10640 20195 10712
rect 15925 6640 16025 10640
rect 20025 6640 20195 10640
rect 15925 6568 20195 6640
rect 20295 6568 20315 10712
rect 15925 6540 20315 6568
rect 20455 10712 24845 10740
rect 20455 10640 24725 10712
rect 20455 6640 20555 10640
rect 24555 6640 24725 10640
rect 20455 6568 24725 6640
rect 24825 6568 24845 10712
rect 20455 6540 24845 6568
rect -24845 6392 -20455 6420
rect -24845 6320 -20575 6392
rect -24845 2320 -24745 6320
rect -20745 2320 -20575 6320
rect -24845 2248 -20575 2320
rect -20475 2248 -20455 6392
rect -24845 2220 -20455 2248
rect -20315 6392 -15925 6420
rect -20315 6320 -16045 6392
rect -20315 2320 -20215 6320
rect -16215 2320 -16045 6320
rect -20315 2248 -16045 2320
rect -15945 2248 -15925 6392
rect -20315 2220 -15925 2248
rect -15785 6392 -11395 6420
rect -15785 6320 -11515 6392
rect -15785 2320 -15685 6320
rect -11685 2320 -11515 6320
rect -15785 2248 -11515 2320
rect -11415 2248 -11395 6392
rect -15785 2220 -11395 2248
rect -11255 6392 -6865 6420
rect -11255 6320 -6985 6392
rect -11255 2320 -11155 6320
rect -7155 2320 -6985 6320
rect -11255 2248 -6985 2320
rect -6885 2248 -6865 6392
rect -11255 2220 -6865 2248
rect -6725 6392 -2335 6420
rect -6725 6320 -2455 6392
rect -6725 2320 -6625 6320
rect -2625 2320 -2455 6320
rect -6725 2248 -2455 2320
rect -2355 2248 -2335 6392
rect -6725 2220 -2335 2248
rect -2195 6392 2195 6420
rect -2195 6320 2075 6392
rect -2195 2320 -2095 6320
rect 1905 2320 2075 6320
rect -2195 2248 2075 2320
rect 2175 2248 2195 6392
rect -2195 2220 2195 2248
rect 2335 6392 6725 6420
rect 2335 6320 6605 6392
rect 2335 2320 2435 6320
rect 6435 2320 6605 6320
rect 2335 2248 6605 2320
rect 6705 2248 6725 6392
rect 2335 2220 6725 2248
rect 6865 6392 11255 6420
rect 6865 6320 11135 6392
rect 6865 2320 6965 6320
rect 10965 2320 11135 6320
rect 6865 2248 11135 2320
rect 11235 2248 11255 6392
rect 6865 2220 11255 2248
rect 11395 6392 15785 6420
rect 11395 6320 15665 6392
rect 11395 2320 11495 6320
rect 15495 2320 15665 6320
rect 11395 2248 15665 2320
rect 15765 2248 15785 6392
rect 11395 2220 15785 2248
rect 15925 6392 20315 6420
rect 15925 6320 20195 6392
rect 15925 2320 16025 6320
rect 20025 2320 20195 6320
rect 15925 2248 20195 2320
rect 20295 2248 20315 6392
rect 15925 2220 20315 2248
rect 20455 6392 24845 6420
rect 20455 6320 24725 6392
rect 20455 2320 20555 6320
rect 24555 2320 24725 6320
rect 20455 2248 24725 2320
rect 24825 2248 24845 6392
rect 20455 2220 24845 2248
rect -24845 2072 -20455 2100
rect -24845 2000 -20575 2072
rect -24845 -2000 -24745 2000
rect -20745 -2000 -20575 2000
rect -24845 -2072 -20575 -2000
rect -20475 -2072 -20455 2072
rect -24845 -2100 -20455 -2072
rect -20315 2072 -15925 2100
rect -20315 2000 -16045 2072
rect -20315 -2000 -20215 2000
rect -16215 -2000 -16045 2000
rect -20315 -2072 -16045 -2000
rect -15945 -2072 -15925 2072
rect -20315 -2100 -15925 -2072
rect -15785 2072 -11395 2100
rect -15785 2000 -11515 2072
rect -15785 -2000 -15685 2000
rect -11685 -2000 -11515 2000
rect -15785 -2072 -11515 -2000
rect -11415 -2072 -11395 2072
rect -15785 -2100 -11395 -2072
rect -11255 2072 -6865 2100
rect -11255 2000 -6985 2072
rect -11255 -2000 -11155 2000
rect -7155 -2000 -6985 2000
rect -11255 -2072 -6985 -2000
rect -6885 -2072 -6865 2072
rect -11255 -2100 -6865 -2072
rect -6725 2072 -2335 2100
rect -6725 2000 -2455 2072
rect -6725 -2000 -6625 2000
rect -2625 -2000 -2455 2000
rect -6725 -2072 -2455 -2000
rect -2355 -2072 -2335 2072
rect -6725 -2100 -2335 -2072
rect -2195 2072 2195 2100
rect -2195 2000 2075 2072
rect -2195 -2000 -2095 2000
rect 1905 -2000 2075 2000
rect -2195 -2072 2075 -2000
rect 2175 -2072 2195 2072
rect -2195 -2100 2195 -2072
rect 2335 2072 6725 2100
rect 2335 2000 6605 2072
rect 2335 -2000 2435 2000
rect 6435 -2000 6605 2000
rect 2335 -2072 6605 -2000
rect 6705 -2072 6725 2072
rect 2335 -2100 6725 -2072
rect 6865 2072 11255 2100
rect 6865 2000 11135 2072
rect 6865 -2000 6965 2000
rect 10965 -2000 11135 2000
rect 6865 -2072 11135 -2000
rect 11235 -2072 11255 2072
rect 6865 -2100 11255 -2072
rect 11395 2072 15785 2100
rect 11395 2000 15665 2072
rect 11395 -2000 11495 2000
rect 15495 -2000 15665 2000
rect 11395 -2072 15665 -2000
rect 15765 -2072 15785 2072
rect 11395 -2100 15785 -2072
rect 15925 2072 20315 2100
rect 15925 2000 20195 2072
rect 15925 -2000 16025 2000
rect 20025 -2000 20195 2000
rect 15925 -2072 20195 -2000
rect 20295 -2072 20315 2072
rect 15925 -2100 20315 -2072
rect 20455 2072 24845 2100
rect 20455 2000 24725 2072
rect 20455 -2000 20555 2000
rect 24555 -2000 24725 2000
rect 20455 -2072 24725 -2000
rect 24825 -2072 24845 2072
rect 20455 -2100 24845 -2072
rect -24845 -2248 -20455 -2220
rect -24845 -2320 -20575 -2248
rect -24845 -6320 -24745 -2320
rect -20745 -6320 -20575 -2320
rect -24845 -6392 -20575 -6320
rect -20475 -6392 -20455 -2248
rect -24845 -6420 -20455 -6392
rect -20315 -2248 -15925 -2220
rect -20315 -2320 -16045 -2248
rect -20315 -6320 -20215 -2320
rect -16215 -6320 -16045 -2320
rect -20315 -6392 -16045 -6320
rect -15945 -6392 -15925 -2248
rect -20315 -6420 -15925 -6392
rect -15785 -2248 -11395 -2220
rect -15785 -2320 -11515 -2248
rect -15785 -6320 -15685 -2320
rect -11685 -6320 -11515 -2320
rect -15785 -6392 -11515 -6320
rect -11415 -6392 -11395 -2248
rect -15785 -6420 -11395 -6392
rect -11255 -2248 -6865 -2220
rect -11255 -2320 -6985 -2248
rect -11255 -6320 -11155 -2320
rect -7155 -6320 -6985 -2320
rect -11255 -6392 -6985 -6320
rect -6885 -6392 -6865 -2248
rect -11255 -6420 -6865 -6392
rect -6725 -2248 -2335 -2220
rect -6725 -2320 -2455 -2248
rect -6725 -6320 -6625 -2320
rect -2625 -6320 -2455 -2320
rect -6725 -6392 -2455 -6320
rect -2355 -6392 -2335 -2248
rect -6725 -6420 -2335 -6392
rect -2195 -2248 2195 -2220
rect -2195 -2320 2075 -2248
rect -2195 -6320 -2095 -2320
rect 1905 -6320 2075 -2320
rect -2195 -6392 2075 -6320
rect 2175 -6392 2195 -2248
rect -2195 -6420 2195 -6392
rect 2335 -2248 6725 -2220
rect 2335 -2320 6605 -2248
rect 2335 -6320 2435 -2320
rect 6435 -6320 6605 -2320
rect 2335 -6392 6605 -6320
rect 6705 -6392 6725 -2248
rect 2335 -6420 6725 -6392
rect 6865 -2248 11255 -2220
rect 6865 -2320 11135 -2248
rect 6865 -6320 6965 -2320
rect 10965 -6320 11135 -2320
rect 6865 -6392 11135 -6320
rect 11235 -6392 11255 -2248
rect 6865 -6420 11255 -6392
rect 11395 -2248 15785 -2220
rect 11395 -2320 15665 -2248
rect 11395 -6320 11495 -2320
rect 15495 -6320 15665 -2320
rect 11395 -6392 15665 -6320
rect 15765 -6392 15785 -2248
rect 11395 -6420 15785 -6392
rect 15925 -2248 20315 -2220
rect 15925 -2320 20195 -2248
rect 15925 -6320 16025 -2320
rect 20025 -6320 20195 -2320
rect 15925 -6392 20195 -6320
rect 20295 -6392 20315 -2248
rect 15925 -6420 20315 -6392
rect 20455 -2248 24845 -2220
rect 20455 -2320 24725 -2248
rect 20455 -6320 20555 -2320
rect 24555 -6320 24725 -2320
rect 20455 -6392 24725 -6320
rect 24825 -6392 24845 -2248
rect 20455 -6420 24845 -6392
rect -24845 -6568 -20455 -6540
rect -24845 -6640 -20575 -6568
rect -24845 -10640 -24745 -6640
rect -20745 -10640 -20575 -6640
rect -24845 -10712 -20575 -10640
rect -20475 -10712 -20455 -6568
rect -24845 -10740 -20455 -10712
rect -20315 -6568 -15925 -6540
rect -20315 -6640 -16045 -6568
rect -20315 -10640 -20215 -6640
rect -16215 -10640 -16045 -6640
rect -20315 -10712 -16045 -10640
rect -15945 -10712 -15925 -6568
rect -20315 -10740 -15925 -10712
rect -15785 -6568 -11395 -6540
rect -15785 -6640 -11515 -6568
rect -15785 -10640 -15685 -6640
rect -11685 -10640 -11515 -6640
rect -15785 -10712 -11515 -10640
rect -11415 -10712 -11395 -6568
rect -15785 -10740 -11395 -10712
rect -11255 -6568 -6865 -6540
rect -11255 -6640 -6985 -6568
rect -11255 -10640 -11155 -6640
rect -7155 -10640 -6985 -6640
rect -11255 -10712 -6985 -10640
rect -6885 -10712 -6865 -6568
rect -11255 -10740 -6865 -10712
rect -6725 -6568 -2335 -6540
rect -6725 -6640 -2455 -6568
rect -6725 -10640 -6625 -6640
rect -2625 -10640 -2455 -6640
rect -6725 -10712 -2455 -10640
rect -2355 -10712 -2335 -6568
rect -6725 -10740 -2335 -10712
rect -2195 -6568 2195 -6540
rect -2195 -6640 2075 -6568
rect -2195 -10640 -2095 -6640
rect 1905 -10640 2075 -6640
rect -2195 -10712 2075 -10640
rect 2175 -10712 2195 -6568
rect -2195 -10740 2195 -10712
rect 2335 -6568 6725 -6540
rect 2335 -6640 6605 -6568
rect 2335 -10640 2435 -6640
rect 6435 -10640 6605 -6640
rect 2335 -10712 6605 -10640
rect 6705 -10712 6725 -6568
rect 2335 -10740 6725 -10712
rect 6865 -6568 11255 -6540
rect 6865 -6640 11135 -6568
rect 6865 -10640 6965 -6640
rect 10965 -10640 11135 -6640
rect 6865 -10712 11135 -10640
rect 11235 -10712 11255 -6568
rect 6865 -10740 11255 -10712
rect 11395 -6568 15785 -6540
rect 11395 -6640 15665 -6568
rect 11395 -10640 11495 -6640
rect 15495 -10640 15665 -6640
rect 11395 -10712 15665 -10640
rect 15765 -10712 15785 -6568
rect 11395 -10740 15785 -10712
rect 15925 -6568 20315 -6540
rect 15925 -6640 20195 -6568
rect 15925 -10640 16025 -6640
rect 20025 -10640 20195 -6640
rect 15925 -10712 20195 -10640
rect 20295 -10712 20315 -6568
rect 15925 -10740 20315 -10712
rect 20455 -6568 24845 -6540
rect 20455 -6640 24725 -6568
rect 20455 -10640 20555 -6640
rect 24555 -10640 24725 -6640
rect 20455 -10712 24725 -10640
rect 24825 -10712 24845 -6568
rect 20455 -10740 24845 -10712
rect -24845 -10888 -20455 -10860
rect -24845 -10960 -20575 -10888
rect -24845 -14960 -24745 -10960
rect -20745 -14960 -20575 -10960
rect -24845 -15032 -20575 -14960
rect -20475 -15032 -20455 -10888
rect -24845 -15060 -20455 -15032
rect -20315 -10888 -15925 -10860
rect -20315 -10960 -16045 -10888
rect -20315 -14960 -20215 -10960
rect -16215 -14960 -16045 -10960
rect -20315 -15032 -16045 -14960
rect -15945 -15032 -15925 -10888
rect -20315 -15060 -15925 -15032
rect -15785 -10888 -11395 -10860
rect -15785 -10960 -11515 -10888
rect -15785 -14960 -15685 -10960
rect -11685 -14960 -11515 -10960
rect -15785 -15032 -11515 -14960
rect -11415 -15032 -11395 -10888
rect -15785 -15060 -11395 -15032
rect -11255 -10888 -6865 -10860
rect -11255 -10960 -6985 -10888
rect -11255 -14960 -11155 -10960
rect -7155 -14960 -6985 -10960
rect -11255 -15032 -6985 -14960
rect -6885 -15032 -6865 -10888
rect -11255 -15060 -6865 -15032
rect -6725 -10888 -2335 -10860
rect -6725 -10960 -2455 -10888
rect -6725 -14960 -6625 -10960
rect -2625 -14960 -2455 -10960
rect -6725 -15032 -2455 -14960
rect -2355 -15032 -2335 -10888
rect -6725 -15060 -2335 -15032
rect -2195 -10888 2195 -10860
rect -2195 -10960 2075 -10888
rect -2195 -14960 -2095 -10960
rect 1905 -14960 2075 -10960
rect -2195 -15032 2075 -14960
rect 2175 -15032 2195 -10888
rect -2195 -15060 2195 -15032
rect 2335 -10888 6725 -10860
rect 2335 -10960 6605 -10888
rect 2335 -14960 2435 -10960
rect 6435 -14960 6605 -10960
rect 2335 -15032 6605 -14960
rect 6705 -15032 6725 -10888
rect 2335 -15060 6725 -15032
rect 6865 -10888 11255 -10860
rect 6865 -10960 11135 -10888
rect 6865 -14960 6965 -10960
rect 10965 -14960 11135 -10960
rect 6865 -15032 11135 -14960
rect 11235 -15032 11255 -10888
rect 6865 -15060 11255 -15032
rect 11395 -10888 15785 -10860
rect 11395 -10960 15665 -10888
rect 11395 -14960 11495 -10960
rect 15495 -14960 15665 -10960
rect 11395 -15032 15665 -14960
rect 15765 -15032 15785 -10888
rect 11395 -15060 15785 -15032
rect 15925 -10888 20315 -10860
rect 15925 -10960 20195 -10888
rect 15925 -14960 16025 -10960
rect 20025 -14960 20195 -10960
rect 15925 -15032 20195 -14960
rect 20295 -15032 20315 -10888
rect 15925 -15060 20315 -15032
rect 20455 -10888 24845 -10860
rect 20455 -10960 24725 -10888
rect 20455 -14960 20555 -10960
rect 24555 -14960 24725 -10960
rect 20455 -15032 24725 -14960
rect 24825 -15032 24845 -10888
rect 20455 -15060 24845 -15032
rect -24845 -15208 -20455 -15180
rect -24845 -15280 -20575 -15208
rect -24845 -19280 -24745 -15280
rect -20745 -19280 -20575 -15280
rect -24845 -19352 -20575 -19280
rect -20475 -19352 -20455 -15208
rect -24845 -19380 -20455 -19352
rect -20315 -15208 -15925 -15180
rect -20315 -15280 -16045 -15208
rect -20315 -19280 -20215 -15280
rect -16215 -19280 -16045 -15280
rect -20315 -19352 -16045 -19280
rect -15945 -19352 -15925 -15208
rect -20315 -19380 -15925 -19352
rect -15785 -15208 -11395 -15180
rect -15785 -15280 -11515 -15208
rect -15785 -19280 -15685 -15280
rect -11685 -19280 -11515 -15280
rect -15785 -19352 -11515 -19280
rect -11415 -19352 -11395 -15208
rect -15785 -19380 -11395 -19352
rect -11255 -15208 -6865 -15180
rect -11255 -15280 -6985 -15208
rect -11255 -19280 -11155 -15280
rect -7155 -19280 -6985 -15280
rect -11255 -19352 -6985 -19280
rect -6885 -19352 -6865 -15208
rect -11255 -19380 -6865 -19352
rect -6725 -15208 -2335 -15180
rect -6725 -15280 -2455 -15208
rect -6725 -19280 -6625 -15280
rect -2625 -19280 -2455 -15280
rect -6725 -19352 -2455 -19280
rect -2355 -19352 -2335 -15208
rect -6725 -19380 -2335 -19352
rect -2195 -15208 2195 -15180
rect -2195 -15280 2075 -15208
rect -2195 -19280 -2095 -15280
rect 1905 -19280 2075 -15280
rect -2195 -19352 2075 -19280
rect 2175 -19352 2195 -15208
rect -2195 -19380 2195 -19352
rect 2335 -15208 6725 -15180
rect 2335 -15280 6605 -15208
rect 2335 -19280 2435 -15280
rect 6435 -19280 6605 -15280
rect 2335 -19352 6605 -19280
rect 6705 -19352 6725 -15208
rect 2335 -19380 6725 -19352
rect 6865 -15208 11255 -15180
rect 6865 -15280 11135 -15208
rect 6865 -19280 6965 -15280
rect 10965 -19280 11135 -15280
rect 6865 -19352 11135 -19280
rect 11235 -19352 11255 -15208
rect 6865 -19380 11255 -19352
rect 11395 -15208 15785 -15180
rect 11395 -15280 15665 -15208
rect 11395 -19280 11495 -15280
rect 15495 -19280 15665 -15280
rect 11395 -19352 15665 -19280
rect 15765 -19352 15785 -15208
rect 11395 -19380 15785 -19352
rect 15925 -15208 20315 -15180
rect 15925 -15280 20195 -15208
rect 15925 -19280 16025 -15280
rect 20025 -19280 20195 -15280
rect 15925 -19352 20195 -19280
rect 20295 -19352 20315 -15208
rect 15925 -19380 20315 -19352
rect 20455 -15208 24845 -15180
rect 20455 -15280 24725 -15208
rect 20455 -19280 20555 -15280
rect 24555 -19280 24725 -15280
rect 20455 -19352 24725 -19280
rect 24825 -19352 24845 -15208
rect 20455 -19380 24845 -19352
rect -24845 -19528 -20455 -19500
rect -24845 -19600 -20575 -19528
rect -24845 -23600 -24745 -19600
rect -20745 -23600 -20575 -19600
rect -24845 -23672 -20575 -23600
rect -20475 -23672 -20455 -19528
rect -24845 -23700 -20455 -23672
rect -20315 -19528 -15925 -19500
rect -20315 -19600 -16045 -19528
rect -20315 -23600 -20215 -19600
rect -16215 -23600 -16045 -19600
rect -20315 -23672 -16045 -23600
rect -15945 -23672 -15925 -19528
rect -20315 -23700 -15925 -23672
rect -15785 -19528 -11395 -19500
rect -15785 -19600 -11515 -19528
rect -15785 -23600 -15685 -19600
rect -11685 -23600 -11515 -19600
rect -15785 -23672 -11515 -23600
rect -11415 -23672 -11395 -19528
rect -15785 -23700 -11395 -23672
rect -11255 -19528 -6865 -19500
rect -11255 -19600 -6985 -19528
rect -11255 -23600 -11155 -19600
rect -7155 -23600 -6985 -19600
rect -11255 -23672 -6985 -23600
rect -6885 -23672 -6865 -19528
rect -11255 -23700 -6865 -23672
rect -6725 -19528 -2335 -19500
rect -6725 -19600 -2455 -19528
rect -6725 -23600 -6625 -19600
rect -2625 -23600 -2455 -19600
rect -6725 -23672 -2455 -23600
rect -2355 -23672 -2335 -19528
rect -6725 -23700 -2335 -23672
rect -2195 -19528 2195 -19500
rect -2195 -19600 2075 -19528
rect -2195 -23600 -2095 -19600
rect 1905 -23600 2075 -19600
rect -2195 -23672 2075 -23600
rect 2175 -23672 2195 -19528
rect -2195 -23700 2195 -23672
rect 2335 -19528 6725 -19500
rect 2335 -19600 6605 -19528
rect 2335 -23600 2435 -19600
rect 6435 -23600 6605 -19600
rect 2335 -23672 6605 -23600
rect 6705 -23672 6725 -19528
rect 2335 -23700 6725 -23672
rect 6865 -19528 11255 -19500
rect 6865 -19600 11135 -19528
rect 6865 -23600 6965 -19600
rect 10965 -23600 11135 -19600
rect 6865 -23672 11135 -23600
rect 11235 -23672 11255 -19528
rect 6865 -23700 11255 -23672
rect 11395 -19528 15785 -19500
rect 11395 -19600 15665 -19528
rect 11395 -23600 11495 -19600
rect 15495 -23600 15665 -19600
rect 11395 -23672 15665 -23600
rect 15765 -23672 15785 -19528
rect 11395 -23700 15785 -23672
rect 15925 -19528 20315 -19500
rect 15925 -19600 20195 -19528
rect 15925 -23600 16025 -19600
rect 20025 -23600 20195 -19600
rect 15925 -23672 20195 -23600
rect 20295 -23672 20315 -19528
rect 15925 -23700 20315 -23672
rect 20455 -19528 24845 -19500
rect 20455 -19600 24725 -19528
rect 20455 -23600 20555 -19600
rect 24555 -23600 24725 -19600
rect 20455 -23672 24725 -23600
rect 24825 -23672 24845 -19528
rect 20455 -23700 24845 -23672
rect -24845 -23848 -20455 -23820
rect -24845 -23920 -20575 -23848
rect -24845 -27920 -24745 -23920
rect -20745 -27920 -20575 -23920
rect -24845 -27992 -20575 -27920
rect -20475 -27992 -20455 -23848
rect -24845 -28020 -20455 -27992
rect -20315 -23848 -15925 -23820
rect -20315 -23920 -16045 -23848
rect -20315 -27920 -20215 -23920
rect -16215 -27920 -16045 -23920
rect -20315 -27992 -16045 -27920
rect -15945 -27992 -15925 -23848
rect -20315 -28020 -15925 -27992
rect -15785 -23848 -11395 -23820
rect -15785 -23920 -11515 -23848
rect -15785 -27920 -15685 -23920
rect -11685 -27920 -11515 -23920
rect -15785 -27992 -11515 -27920
rect -11415 -27992 -11395 -23848
rect -15785 -28020 -11395 -27992
rect -11255 -23848 -6865 -23820
rect -11255 -23920 -6985 -23848
rect -11255 -27920 -11155 -23920
rect -7155 -27920 -6985 -23920
rect -11255 -27992 -6985 -27920
rect -6885 -27992 -6865 -23848
rect -11255 -28020 -6865 -27992
rect -6725 -23848 -2335 -23820
rect -6725 -23920 -2455 -23848
rect -6725 -27920 -6625 -23920
rect -2625 -27920 -2455 -23920
rect -6725 -27992 -2455 -27920
rect -2355 -27992 -2335 -23848
rect -6725 -28020 -2335 -27992
rect -2195 -23848 2195 -23820
rect -2195 -23920 2075 -23848
rect -2195 -27920 -2095 -23920
rect 1905 -27920 2075 -23920
rect -2195 -27992 2075 -27920
rect 2175 -27992 2195 -23848
rect -2195 -28020 2195 -27992
rect 2335 -23848 6725 -23820
rect 2335 -23920 6605 -23848
rect 2335 -27920 2435 -23920
rect 6435 -27920 6605 -23920
rect 2335 -27992 6605 -27920
rect 6705 -27992 6725 -23848
rect 2335 -28020 6725 -27992
rect 6865 -23848 11255 -23820
rect 6865 -23920 11135 -23848
rect 6865 -27920 6965 -23920
rect 10965 -27920 11135 -23920
rect 6865 -27992 11135 -27920
rect 11235 -27992 11255 -23848
rect 6865 -28020 11255 -27992
rect 11395 -23848 15785 -23820
rect 11395 -23920 15665 -23848
rect 11395 -27920 11495 -23920
rect 15495 -27920 15665 -23920
rect 11395 -27992 15665 -27920
rect 15765 -27992 15785 -23848
rect 11395 -28020 15785 -27992
rect 15925 -23848 20315 -23820
rect 15925 -23920 20195 -23848
rect 15925 -27920 16025 -23920
rect 20025 -27920 20195 -23920
rect 15925 -27992 20195 -27920
rect 20295 -27992 20315 -23848
rect 15925 -28020 20315 -27992
rect 20455 -23848 24845 -23820
rect 20455 -23920 24725 -23848
rect 20455 -27920 20555 -23920
rect 24555 -27920 24725 -23920
rect 20455 -27992 24725 -27920
rect 24825 -27992 24845 -23848
rect 20455 -28020 24845 -27992
rect -24845 -28168 -20455 -28140
rect -24845 -28240 -20575 -28168
rect -24845 -32240 -24745 -28240
rect -20745 -32240 -20575 -28240
rect -24845 -32312 -20575 -32240
rect -20475 -32312 -20455 -28168
rect -24845 -32340 -20455 -32312
rect -20315 -28168 -15925 -28140
rect -20315 -28240 -16045 -28168
rect -20315 -32240 -20215 -28240
rect -16215 -32240 -16045 -28240
rect -20315 -32312 -16045 -32240
rect -15945 -32312 -15925 -28168
rect -20315 -32340 -15925 -32312
rect -15785 -28168 -11395 -28140
rect -15785 -28240 -11515 -28168
rect -15785 -32240 -15685 -28240
rect -11685 -32240 -11515 -28240
rect -15785 -32312 -11515 -32240
rect -11415 -32312 -11395 -28168
rect -15785 -32340 -11395 -32312
rect -11255 -28168 -6865 -28140
rect -11255 -28240 -6985 -28168
rect -11255 -32240 -11155 -28240
rect -7155 -32240 -6985 -28240
rect -11255 -32312 -6985 -32240
rect -6885 -32312 -6865 -28168
rect -11255 -32340 -6865 -32312
rect -6725 -28168 -2335 -28140
rect -6725 -28240 -2455 -28168
rect -6725 -32240 -6625 -28240
rect -2625 -32240 -2455 -28240
rect -6725 -32312 -2455 -32240
rect -2355 -32312 -2335 -28168
rect -6725 -32340 -2335 -32312
rect -2195 -28168 2195 -28140
rect -2195 -28240 2075 -28168
rect -2195 -32240 -2095 -28240
rect 1905 -32240 2075 -28240
rect -2195 -32312 2075 -32240
rect 2175 -32312 2195 -28168
rect -2195 -32340 2195 -32312
rect 2335 -28168 6725 -28140
rect 2335 -28240 6605 -28168
rect 2335 -32240 2435 -28240
rect 6435 -32240 6605 -28240
rect 2335 -32312 6605 -32240
rect 6705 -32312 6725 -28168
rect 2335 -32340 6725 -32312
rect 6865 -28168 11255 -28140
rect 6865 -28240 11135 -28168
rect 6865 -32240 6965 -28240
rect 10965 -32240 11135 -28240
rect 6865 -32312 11135 -32240
rect 11235 -32312 11255 -28168
rect 6865 -32340 11255 -32312
rect 11395 -28168 15785 -28140
rect 11395 -28240 15665 -28168
rect 11395 -32240 11495 -28240
rect 15495 -32240 15665 -28240
rect 11395 -32312 15665 -32240
rect 15765 -32312 15785 -28168
rect 11395 -32340 15785 -32312
rect 15925 -28168 20315 -28140
rect 15925 -28240 20195 -28168
rect 15925 -32240 16025 -28240
rect 20025 -32240 20195 -28240
rect 15925 -32312 20195 -32240
rect 20295 -32312 20315 -28168
rect 15925 -32340 20315 -32312
rect 20455 -28168 24845 -28140
rect 20455 -28240 24725 -28168
rect 20455 -32240 20555 -28240
rect 24555 -32240 24725 -28240
rect 20455 -32312 24725 -32240
rect 24825 -32312 24845 -28168
rect 20455 -32340 24845 -32312
<< viatp >>
rect -20575 28168 -20475 32312
rect -16045 28168 -15945 32312
rect -11515 28168 -11415 32312
rect -6985 28168 -6885 32312
rect -2455 28168 -2355 32312
rect 2075 28168 2175 32312
rect 6605 28168 6705 32312
rect 11135 28168 11235 32312
rect 15665 28168 15765 32312
rect 20195 28168 20295 32312
rect 24725 28168 24825 32312
rect -20575 23848 -20475 27992
rect -16045 23848 -15945 27992
rect -11515 23848 -11415 27992
rect -6985 23848 -6885 27992
rect -2455 23848 -2355 27992
rect 2075 23848 2175 27992
rect 6605 23848 6705 27992
rect 11135 23848 11235 27992
rect 15665 23848 15765 27992
rect 20195 23848 20295 27992
rect 24725 23848 24825 27992
rect -20575 19528 -20475 23672
rect -16045 19528 -15945 23672
rect -11515 19528 -11415 23672
rect -6985 19528 -6885 23672
rect -2455 19528 -2355 23672
rect 2075 19528 2175 23672
rect 6605 19528 6705 23672
rect 11135 19528 11235 23672
rect 15665 19528 15765 23672
rect 20195 19528 20295 23672
rect 24725 19528 24825 23672
rect -20575 15208 -20475 19352
rect -16045 15208 -15945 19352
rect -11515 15208 -11415 19352
rect -6985 15208 -6885 19352
rect -2455 15208 -2355 19352
rect 2075 15208 2175 19352
rect 6605 15208 6705 19352
rect 11135 15208 11235 19352
rect 15665 15208 15765 19352
rect 20195 15208 20295 19352
rect 24725 15208 24825 19352
rect -20575 10888 -20475 15032
rect -16045 10888 -15945 15032
rect -11515 10888 -11415 15032
rect -6985 10888 -6885 15032
rect -2455 10888 -2355 15032
rect 2075 10888 2175 15032
rect 6605 10888 6705 15032
rect 11135 10888 11235 15032
rect 15665 10888 15765 15032
rect 20195 10888 20295 15032
rect 24725 10888 24825 15032
rect -20575 6568 -20475 10712
rect -16045 6568 -15945 10712
rect -11515 6568 -11415 10712
rect -6985 6568 -6885 10712
rect -2455 6568 -2355 10712
rect 2075 6568 2175 10712
rect 6605 6568 6705 10712
rect 11135 6568 11235 10712
rect 15665 6568 15765 10712
rect 20195 6568 20295 10712
rect 24725 6568 24825 10712
rect -20575 2248 -20475 6392
rect -16045 2248 -15945 6392
rect -11515 2248 -11415 6392
rect -6985 2248 -6885 6392
rect -2455 2248 -2355 6392
rect 2075 2248 2175 6392
rect 6605 2248 6705 6392
rect 11135 2248 11235 6392
rect 15665 2248 15765 6392
rect 20195 2248 20295 6392
rect 24725 2248 24825 6392
rect -20575 -2072 -20475 2072
rect -16045 -2072 -15945 2072
rect -11515 -2072 -11415 2072
rect -6985 -2072 -6885 2072
rect -2455 -2072 -2355 2072
rect 2075 -2072 2175 2072
rect 6605 -2072 6705 2072
rect 11135 -2072 11235 2072
rect 15665 -2072 15765 2072
rect 20195 -2072 20295 2072
rect 24725 -2072 24825 2072
rect -20575 -6392 -20475 -2248
rect -16045 -6392 -15945 -2248
rect -11515 -6392 -11415 -2248
rect -6985 -6392 -6885 -2248
rect -2455 -6392 -2355 -2248
rect 2075 -6392 2175 -2248
rect 6605 -6392 6705 -2248
rect 11135 -6392 11235 -2248
rect 15665 -6392 15765 -2248
rect 20195 -6392 20295 -2248
rect 24725 -6392 24825 -2248
rect -20575 -10712 -20475 -6568
rect -16045 -10712 -15945 -6568
rect -11515 -10712 -11415 -6568
rect -6985 -10712 -6885 -6568
rect -2455 -10712 -2355 -6568
rect 2075 -10712 2175 -6568
rect 6605 -10712 6705 -6568
rect 11135 -10712 11235 -6568
rect 15665 -10712 15765 -6568
rect 20195 -10712 20295 -6568
rect 24725 -10712 24825 -6568
rect -20575 -15032 -20475 -10888
rect -16045 -15032 -15945 -10888
rect -11515 -15032 -11415 -10888
rect -6985 -15032 -6885 -10888
rect -2455 -15032 -2355 -10888
rect 2075 -15032 2175 -10888
rect 6605 -15032 6705 -10888
rect 11135 -15032 11235 -10888
rect 15665 -15032 15765 -10888
rect 20195 -15032 20295 -10888
rect 24725 -15032 24825 -10888
rect -20575 -19352 -20475 -15208
rect -16045 -19352 -15945 -15208
rect -11515 -19352 -11415 -15208
rect -6985 -19352 -6885 -15208
rect -2455 -19352 -2355 -15208
rect 2075 -19352 2175 -15208
rect 6605 -19352 6705 -15208
rect 11135 -19352 11235 -15208
rect 15665 -19352 15765 -15208
rect 20195 -19352 20295 -15208
rect 24725 -19352 24825 -15208
rect -20575 -23672 -20475 -19528
rect -16045 -23672 -15945 -19528
rect -11515 -23672 -11415 -19528
rect -6985 -23672 -6885 -19528
rect -2455 -23672 -2355 -19528
rect 2075 -23672 2175 -19528
rect 6605 -23672 6705 -19528
rect 11135 -23672 11235 -19528
rect 15665 -23672 15765 -19528
rect 20195 -23672 20295 -19528
rect 24725 -23672 24825 -19528
rect -20575 -27992 -20475 -23848
rect -16045 -27992 -15945 -23848
rect -11515 -27992 -11415 -23848
rect -6985 -27992 -6885 -23848
rect -2455 -27992 -2355 -23848
rect 2075 -27992 2175 -23848
rect 6605 -27992 6705 -23848
rect 11135 -27992 11235 -23848
rect 15665 -27992 15765 -23848
rect 20195 -27992 20295 -23848
rect 24725 -27992 24825 -23848
rect -20575 -32312 -20475 -28168
rect -16045 -32312 -15945 -28168
rect -11515 -32312 -11415 -28168
rect -6985 -32312 -6885 -28168
rect -2455 -32312 -2355 -28168
rect 2075 -32312 2175 -28168
rect 6605 -32312 6705 -28168
rect 11135 -32312 11235 -28168
rect 15665 -32312 15765 -28168
rect 20195 -32312 20295 -28168
rect 24725 -32312 24825 -28168
<< metaltp >>
rect -22815 32210 -22675 32400
rect -20595 32312 -20455 32400
rect -22815 27890 -22675 28270
rect -20595 28168 -20575 32312
rect -20475 28168 -20455 32312
rect -18285 32210 -18145 32400
rect -16065 32312 -15925 32400
rect -20595 27992 -20455 28168
rect -22815 23570 -22675 23950
rect -20595 23848 -20575 27992
rect -20475 23848 -20455 27992
rect -18285 27890 -18145 28270
rect -16065 28168 -16045 32312
rect -15945 28168 -15925 32312
rect -13755 32210 -13615 32400
rect -11535 32312 -11395 32400
rect -16065 27992 -15925 28168
rect -20595 23672 -20455 23848
rect -22815 19250 -22675 19630
rect -20595 19528 -20575 23672
rect -20475 19528 -20455 23672
rect -18285 23570 -18145 23950
rect -16065 23848 -16045 27992
rect -15945 23848 -15925 27992
rect -13755 27890 -13615 28270
rect -11535 28168 -11515 32312
rect -11415 28168 -11395 32312
rect -9225 32210 -9085 32400
rect -7005 32312 -6865 32400
rect -11535 27992 -11395 28168
rect -16065 23672 -15925 23848
rect -20595 19352 -20455 19528
rect -22815 14930 -22675 15310
rect -20595 15208 -20575 19352
rect -20475 15208 -20455 19352
rect -18285 19250 -18145 19630
rect -16065 19528 -16045 23672
rect -15945 19528 -15925 23672
rect -13755 23570 -13615 23950
rect -11535 23848 -11515 27992
rect -11415 23848 -11395 27992
rect -9225 27890 -9085 28270
rect -7005 28168 -6985 32312
rect -6885 28168 -6865 32312
rect -4695 32210 -4555 32400
rect -2475 32312 -2335 32400
rect -7005 27992 -6865 28168
rect -11535 23672 -11395 23848
rect -16065 19352 -15925 19528
rect -20595 15032 -20455 15208
rect -22815 10610 -22675 10990
rect -20595 10888 -20575 15032
rect -20475 10888 -20455 15032
rect -18285 14930 -18145 15310
rect -16065 15208 -16045 19352
rect -15945 15208 -15925 19352
rect -13755 19250 -13615 19630
rect -11535 19528 -11515 23672
rect -11415 19528 -11395 23672
rect -9225 23570 -9085 23950
rect -7005 23848 -6985 27992
rect -6885 23848 -6865 27992
rect -4695 27890 -4555 28270
rect -2475 28168 -2455 32312
rect -2355 28168 -2335 32312
rect -165 32210 -25 32400
rect 2055 32312 2195 32400
rect -2475 27992 -2335 28168
rect -7005 23672 -6865 23848
rect -11535 19352 -11395 19528
rect -16065 15032 -15925 15208
rect -20595 10712 -20455 10888
rect -22815 6290 -22675 6670
rect -20595 6568 -20575 10712
rect -20475 6568 -20455 10712
rect -18285 10610 -18145 10990
rect -16065 10888 -16045 15032
rect -15945 10888 -15925 15032
rect -13755 14930 -13615 15310
rect -11535 15208 -11515 19352
rect -11415 15208 -11395 19352
rect -9225 19250 -9085 19630
rect -7005 19528 -6985 23672
rect -6885 19528 -6865 23672
rect -4695 23570 -4555 23950
rect -2475 23848 -2455 27992
rect -2355 23848 -2335 27992
rect -165 27890 -25 28270
rect 2055 28168 2075 32312
rect 2175 28168 2195 32312
rect 4365 32210 4505 32400
rect 6585 32312 6725 32400
rect 2055 27992 2195 28168
rect -2475 23672 -2335 23848
rect -7005 19352 -6865 19528
rect -11535 15032 -11395 15208
rect -16065 10712 -15925 10888
rect -20595 6392 -20455 6568
rect -22815 1970 -22675 2350
rect -20595 2248 -20575 6392
rect -20475 2248 -20455 6392
rect -18285 6290 -18145 6670
rect -16065 6568 -16045 10712
rect -15945 6568 -15925 10712
rect -13755 10610 -13615 10990
rect -11535 10888 -11515 15032
rect -11415 10888 -11395 15032
rect -9225 14930 -9085 15310
rect -7005 15208 -6985 19352
rect -6885 15208 -6865 19352
rect -4695 19250 -4555 19630
rect -2475 19528 -2455 23672
rect -2355 19528 -2335 23672
rect -165 23570 -25 23950
rect 2055 23848 2075 27992
rect 2175 23848 2195 27992
rect 4365 27890 4505 28270
rect 6585 28168 6605 32312
rect 6705 28168 6725 32312
rect 8895 32210 9035 32400
rect 11115 32312 11255 32400
rect 6585 27992 6725 28168
rect 2055 23672 2195 23848
rect -2475 19352 -2335 19528
rect -7005 15032 -6865 15208
rect -11535 10712 -11395 10888
rect -16065 6392 -15925 6568
rect -20595 2072 -20455 2248
rect -22815 -2350 -22675 -1970
rect -20595 -2072 -20575 2072
rect -20475 -2072 -20455 2072
rect -18285 1970 -18145 2350
rect -16065 2248 -16045 6392
rect -15945 2248 -15925 6392
rect -13755 6290 -13615 6670
rect -11535 6568 -11515 10712
rect -11415 6568 -11395 10712
rect -9225 10610 -9085 10990
rect -7005 10888 -6985 15032
rect -6885 10888 -6865 15032
rect -4695 14930 -4555 15310
rect -2475 15208 -2455 19352
rect -2355 15208 -2335 19352
rect -165 19250 -25 19630
rect 2055 19528 2075 23672
rect 2175 19528 2195 23672
rect 4365 23570 4505 23950
rect 6585 23848 6605 27992
rect 6705 23848 6725 27992
rect 8895 27890 9035 28270
rect 11115 28168 11135 32312
rect 11235 28168 11255 32312
rect 13425 32210 13565 32400
rect 15645 32312 15785 32400
rect 11115 27992 11255 28168
rect 6585 23672 6725 23848
rect 2055 19352 2195 19528
rect -2475 15032 -2335 15208
rect -7005 10712 -6865 10888
rect -11535 6392 -11395 6568
rect -16065 2072 -15925 2248
rect -20595 -2248 -20455 -2072
rect -22815 -6670 -22675 -6290
rect -20595 -6392 -20575 -2248
rect -20475 -6392 -20455 -2248
rect -18285 -2350 -18145 -1970
rect -16065 -2072 -16045 2072
rect -15945 -2072 -15925 2072
rect -13755 1970 -13615 2350
rect -11535 2248 -11515 6392
rect -11415 2248 -11395 6392
rect -9225 6290 -9085 6670
rect -7005 6568 -6985 10712
rect -6885 6568 -6865 10712
rect -4695 10610 -4555 10990
rect -2475 10888 -2455 15032
rect -2355 10888 -2335 15032
rect -165 14930 -25 15310
rect 2055 15208 2075 19352
rect 2175 15208 2195 19352
rect 4365 19250 4505 19630
rect 6585 19528 6605 23672
rect 6705 19528 6725 23672
rect 8895 23570 9035 23950
rect 11115 23848 11135 27992
rect 11235 23848 11255 27992
rect 13425 27890 13565 28270
rect 15645 28168 15665 32312
rect 15765 28168 15785 32312
rect 17955 32210 18095 32400
rect 20175 32312 20315 32400
rect 15645 27992 15785 28168
rect 11115 23672 11255 23848
rect 6585 19352 6725 19528
rect 2055 15032 2195 15208
rect -2475 10712 -2335 10888
rect -7005 6392 -6865 6568
rect -11535 2072 -11395 2248
rect -16065 -2248 -15925 -2072
rect -20595 -6568 -20455 -6392
rect -22815 -10990 -22675 -10610
rect -20595 -10712 -20575 -6568
rect -20475 -10712 -20455 -6568
rect -18285 -6670 -18145 -6290
rect -16065 -6392 -16045 -2248
rect -15945 -6392 -15925 -2248
rect -13755 -2350 -13615 -1970
rect -11535 -2072 -11515 2072
rect -11415 -2072 -11395 2072
rect -9225 1970 -9085 2350
rect -7005 2248 -6985 6392
rect -6885 2248 -6865 6392
rect -4695 6290 -4555 6670
rect -2475 6568 -2455 10712
rect -2355 6568 -2335 10712
rect -165 10610 -25 10990
rect 2055 10888 2075 15032
rect 2175 10888 2195 15032
rect 4365 14930 4505 15310
rect 6585 15208 6605 19352
rect 6705 15208 6725 19352
rect 8895 19250 9035 19630
rect 11115 19528 11135 23672
rect 11235 19528 11255 23672
rect 13425 23570 13565 23950
rect 15645 23848 15665 27992
rect 15765 23848 15785 27992
rect 17955 27890 18095 28270
rect 20175 28168 20195 32312
rect 20295 28168 20315 32312
rect 22485 32210 22625 32400
rect 24705 32312 24845 32400
rect 20175 27992 20315 28168
rect 15645 23672 15785 23848
rect 11115 19352 11255 19528
rect 6585 15032 6725 15208
rect 2055 10712 2195 10888
rect -2475 6392 -2335 6568
rect -7005 2072 -6865 2248
rect -11535 -2248 -11395 -2072
rect -16065 -6568 -15925 -6392
rect -20595 -10888 -20455 -10712
rect -22815 -15310 -22675 -14930
rect -20595 -15032 -20575 -10888
rect -20475 -15032 -20455 -10888
rect -18285 -10990 -18145 -10610
rect -16065 -10712 -16045 -6568
rect -15945 -10712 -15925 -6568
rect -13755 -6670 -13615 -6290
rect -11535 -6392 -11515 -2248
rect -11415 -6392 -11395 -2248
rect -9225 -2350 -9085 -1970
rect -7005 -2072 -6985 2072
rect -6885 -2072 -6865 2072
rect -4695 1970 -4555 2350
rect -2475 2248 -2455 6392
rect -2355 2248 -2335 6392
rect -165 6290 -25 6670
rect 2055 6568 2075 10712
rect 2175 6568 2195 10712
rect 4365 10610 4505 10990
rect 6585 10888 6605 15032
rect 6705 10888 6725 15032
rect 8895 14930 9035 15310
rect 11115 15208 11135 19352
rect 11235 15208 11255 19352
rect 13425 19250 13565 19630
rect 15645 19528 15665 23672
rect 15765 19528 15785 23672
rect 17955 23570 18095 23950
rect 20175 23848 20195 27992
rect 20295 23848 20315 27992
rect 22485 27890 22625 28270
rect 24705 28168 24725 32312
rect 24825 28168 24845 32312
rect 24705 27992 24845 28168
rect 20175 23672 20315 23848
rect 15645 19352 15785 19528
rect 11115 15032 11255 15208
rect 6585 10712 6725 10888
rect 2055 6392 2195 6568
rect -2475 2072 -2335 2248
rect -7005 -2248 -6865 -2072
rect -11535 -6568 -11395 -6392
rect -16065 -10888 -15925 -10712
rect -20595 -15208 -20455 -15032
rect -22815 -19630 -22675 -19250
rect -20595 -19352 -20575 -15208
rect -20475 -19352 -20455 -15208
rect -18285 -15310 -18145 -14930
rect -16065 -15032 -16045 -10888
rect -15945 -15032 -15925 -10888
rect -13755 -10990 -13615 -10610
rect -11535 -10712 -11515 -6568
rect -11415 -10712 -11395 -6568
rect -9225 -6670 -9085 -6290
rect -7005 -6392 -6985 -2248
rect -6885 -6392 -6865 -2248
rect -4695 -2350 -4555 -1970
rect -2475 -2072 -2455 2072
rect -2355 -2072 -2335 2072
rect -165 1970 -25 2350
rect 2055 2248 2075 6392
rect 2175 2248 2195 6392
rect 4365 6290 4505 6670
rect 6585 6568 6605 10712
rect 6705 6568 6725 10712
rect 8895 10610 9035 10990
rect 11115 10888 11135 15032
rect 11235 10888 11255 15032
rect 13425 14930 13565 15310
rect 15645 15208 15665 19352
rect 15765 15208 15785 19352
rect 17955 19250 18095 19630
rect 20175 19528 20195 23672
rect 20295 19528 20315 23672
rect 22485 23570 22625 23950
rect 24705 23848 24725 27992
rect 24825 23848 24845 27992
rect 24705 23672 24845 23848
rect 20175 19352 20315 19528
rect 15645 15032 15785 15208
rect 11115 10712 11255 10888
rect 6585 6392 6725 6568
rect 2055 2072 2195 2248
rect -2475 -2248 -2335 -2072
rect -7005 -6568 -6865 -6392
rect -11535 -10888 -11395 -10712
rect -16065 -15208 -15925 -15032
rect -20595 -19528 -20455 -19352
rect -22815 -23950 -22675 -23570
rect -20595 -23672 -20575 -19528
rect -20475 -23672 -20455 -19528
rect -18285 -19630 -18145 -19250
rect -16065 -19352 -16045 -15208
rect -15945 -19352 -15925 -15208
rect -13755 -15310 -13615 -14930
rect -11535 -15032 -11515 -10888
rect -11415 -15032 -11395 -10888
rect -9225 -10990 -9085 -10610
rect -7005 -10712 -6985 -6568
rect -6885 -10712 -6865 -6568
rect -4695 -6670 -4555 -6290
rect -2475 -6392 -2455 -2248
rect -2355 -6392 -2335 -2248
rect -165 -2350 -25 -1970
rect 2055 -2072 2075 2072
rect 2175 -2072 2195 2072
rect 4365 1970 4505 2350
rect 6585 2248 6605 6392
rect 6705 2248 6725 6392
rect 8895 6290 9035 6670
rect 11115 6568 11135 10712
rect 11235 6568 11255 10712
rect 13425 10610 13565 10990
rect 15645 10888 15665 15032
rect 15765 10888 15785 15032
rect 17955 14930 18095 15310
rect 20175 15208 20195 19352
rect 20295 15208 20315 19352
rect 22485 19250 22625 19630
rect 24705 19528 24725 23672
rect 24825 19528 24845 23672
rect 24705 19352 24845 19528
rect 20175 15032 20315 15208
rect 15645 10712 15785 10888
rect 11115 6392 11255 6568
rect 6585 2072 6725 2248
rect 2055 -2248 2195 -2072
rect -2475 -6568 -2335 -6392
rect -7005 -10888 -6865 -10712
rect -11535 -15208 -11395 -15032
rect -16065 -19528 -15925 -19352
rect -20595 -23848 -20455 -23672
rect -22815 -28270 -22675 -27890
rect -20595 -27992 -20575 -23848
rect -20475 -27992 -20455 -23848
rect -18285 -23950 -18145 -23570
rect -16065 -23672 -16045 -19528
rect -15945 -23672 -15925 -19528
rect -13755 -19630 -13615 -19250
rect -11535 -19352 -11515 -15208
rect -11415 -19352 -11395 -15208
rect -9225 -15310 -9085 -14930
rect -7005 -15032 -6985 -10888
rect -6885 -15032 -6865 -10888
rect -4695 -10990 -4555 -10610
rect -2475 -10712 -2455 -6568
rect -2355 -10712 -2335 -6568
rect -165 -6670 -25 -6290
rect 2055 -6392 2075 -2248
rect 2175 -6392 2195 -2248
rect 4365 -2350 4505 -1970
rect 6585 -2072 6605 2072
rect 6705 -2072 6725 2072
rect 8895 1970 9035 2350
rect 11115 2248 11135 6392
rect 11235 2248 11255 6392
rect 13425 6290 13565 6670
rect 15645 6568 15665 10712
rect 15765 6568 15785 10712
rect 17955 10610 18095 10990
rect 20175 10888 20195 15032
rect 20295 10888 20315 15032
rect 22485 14930 22625 15310
rect 24705 15208 24725 19352
rect 24825 15208 24845 19352
rect 24705 15032 24845 15208
rect 20175 10712 20315 10888
rect 15645 6392 15785 6568
rect 11115 2072 11255 2248
rect 6585 -2248 6725 -2072
rect 2055 -6568 2195 -6392
rect -2475 -10888 -2335 -10712
rect -7005 -15208 -6865 -15032
rect -11535 -19528 -11395 -19352
rect -16065 -23848 -15925 -23672
rect -20595 -28168 -20455 -27992
rect -22815 -32400 -22675 -32210
rect -20595 -32312 -20575 -28168
rect -20475 -32312 -20455 -28168
rect -18285 -28270 -18145 -27890
rect -16065 -27992 -16045 -23848
rect -15945 -27992 -15925 -23848
rect -13755 -23950 -13615 -23570
rect -11535 -23672 -11515 -19528
rect -11415 -23672 -11395 -19528
rect -9225 -19630 -9085 -19250
rect -7005 -19352 -6985 -15208
rect -6885 -19352 -6865 -15208
rect -4695 -15310 -4555 -14930
rect -2475 -15032 -2455 -10888
rect -2355 -15032 -2335 -10888
rect -165 -10990 -25 -10610
rect 2055 -10712 2075 -6568
rect 2175 -10712 2195 -6568
rect 4365 -6670 4505 -6290
rect 6585 -6392 6605 -2248
rect 6705 -6392 6725 -2248
rect 8895 -2350 9035 -1970
rect 11115 -2072 11135 2072
rect 11235 -2072 11255 2072
rect 13425 1970 13565 2350
rect 15645 2248 15665 6392
rect 15765 2248 15785 6392
rect 17955 6290 18095 6670
rect 20175 6568 20195 10712
rect 20295 6568 20315 10712
rect 22485 10610 22625 10990
rect 24705 10888 24725 15032
rect 24825 10888 24845 15032
rect 24705 10712 24845 10888
rect 20175 6392 20315 6568
rect 15645 2072 15785 2248
rect 11115 -2248 11255 -2072
rect 6585 -6568 6725 -6392
rect 2055 -10888 2195 -10712
rect -2475 -15208 -2335 -15032
rect -7005 -19528 -6865 -19352
rect -11535 -23848 -11395 -23672
rect -16065 -28168 -15925 -27992
rect -20595 -32400 -20455 -32312
rect -18285 -32400 -18145 -32210
rect -16065 -32312 -16045 -28168
rect -15945 -32312 -15925 -28168
rect -13755 -28270 -13615 -27890
rect -11535 -27992 -11515 -23848
rect -11415 -27992 -11395 -23848
rect -9225 -23950 -9085 -23570
rect -7005 -23672 -6985 -19528
rect -6885 -23672 -6865 -19528
rect -4695 -19630 -4555 -19250
rect -2475 -19352 -2455 -15208
rect -2355 -19352 -2335 -15208
rect -165 -15310 -25 -14930
rect 2055 -15032 2075 -10888
rect 2175 -15032 2195 -10888
rect 4365 -10990 4505 -10610
rect 6585 -10712 6605 -6568
rect 6705 -10712 6725 -6568
rect 8895 -6670 9035 -6290
rect 11115 -6392 11135 -2248
rect 11235 -6392 11255 -2248
rect 13425 -2350 13565 -1970
rect 15645 -2072 15665 2072
rect 15765 -2072 15785 2072
rect 17955 1970 18095 2350
rect 20175 2248 20195 6392
rect 20295 2248 20315 6392
rect 22485 6290 22625 6670
rect 24705 6568 24725 10712
rect 24825 6568 24845 10712
rect 24705 6392 24845 6568
rect 20175 2072 20315 2248
rect 15645 -2248 15785 -2072
rect 11115 -6568 11255 -6392
rect 6585 -10888 6725 -10712
rect 2055 -15208 2195 -15032
rect -2475 -19528 -2335 -19352
rect -7005 -23848 -6865 -23672
rect -11535 -28168 -11395 -27992
rect -16065 -32400 -15925 -32312
rect -13755 -32400 -13615 -32210
rect -11535 -32312 -11515 -28168
rect -11415 -32312 -11395 -28168
rect -9225 -28270 -9085 -27890
rect -7005 -27992 -6985 -23848
rect -6885 -27992 -6865 -23848
rect -4695 -23950 -4555 -23570
rect -2475 -23672 -2455 -19528
rect -2355 -23672 -2335 -19528
rect -165 -19630 -25 -19250
rect 2055 -19352 2075 -15208
rect 2175 -19352 2195 -15208
rect 4365 -15310 4505 -14930
rect 6585 -15032 6605 -10888
rect 6705 -15032 6725 -10888
rect 8895 -10990 9035 -10610
rect 11115 -10712 11135 -6568
rect 11235 -10712 11255 -6568
rect 13425 -6670 13565 -6290
rect 15645 -6392 15665 -2248
rect 15765 -6392 15785 -2248
rect 17955 -2350 18095 -1970
rect 20175 -2072 20195 2072
rect 20295 -2072 20315 2072
rect 22485 1970 22625 2350
rect 24705 2248 24725 6392
rect 24825 2248 24845 6392
rect 24705 2072 24845 2248
rect 20175 -2248 20315 -2072
rect 15645 -6568 15785 -6392
rect 11115 -10888 11255 -10712
rect 6585 -15208 6725 -15032
rect 2055 -19528 2195 -19352
rect -2475 -23848 -2335 -23672
rect -7005 -28168 -6865 -27992
rect -11535 -32400 -11395 -32312
rect -9225 -32400 -9085 -32210
rect -7005 -32312 -6985 -28168
rect -6885 -32312 -6865 -28168
rect -4695 -28270 -4555 -27890
rect -2475 -27992 -2455 -23848
rect -2355 -27992 -2335 -23848
rect -165 -23950 -25 -23570
rect 2055 -23672 2075 -19528
rect 2175 -23672 2195 -19528
rect 4365 -19630 4505 -19250
rect 6585 -19352 6605 -15208
rect 6705 -19352 6725 -15208
rect 8895 -15310 9035 -14930
rect 11115 -15032 11135 -10888
rect 11235 -15032 11255 -10888
rect 13425 -10990 13565 -10610
rect 15645 -10712 15665 -6568
rect 15765 -10712 15785 -6568
rect 17955 -6670 18095 -6290
rect 20175 -6392 20195 -2248
rect 20295 -6392 20315 -2248
rect 22485 -2350 22625 -1970
rect 24705 -2072 24725 2072
rect 24825 -2072 24845 2072
rect 24705 -2248 24845 -2072
rect 20175 -6568 20315 -6392
rect 15645 -10888 15785 -10712
rect 11115 -15208 11255 -15032
rect 6585 -19528 6725 -19352
rect 2055 -23848 2195 -23672
rect -2475 -28168 -2335 -27992
rect -7005 -32400 -6865 -32312
rect -4695 -32400 -4555 -32210
rect -2475 -32312 -2455 -28168
rect -2355 -32312 -2335 -28168
rect -165 -28270 -25 -27890
rect 2055 -27992 2075 -23848
rect 2175 -27992 2195 -23848
rect 4365 -23950 4505 -23570
rect 6585 -23672 6605 -19528
rect 6705 -23672 6725 -19528
rect 8895 -19630 9035 -19250
rect 11115 -19352 11135 -15208
rect 11235 -19352 11255 -15208
rect 13425 -15310 13565 -14930
rect 15645 -15032 15665 -10888
rect 15765 -15032 15785 -10888
rect 17955 -10990 18095 -10610
rect 20175 -10712 20195 -6568
rect 20295 -10712 20315 -6568
rect 22485 -6670 22625 -6290
rect 24705 -6392 24725 -2248
rect 24825 -6392 24845 -2248
rect 24705 -6568 24845 -6392
rect 20175 -10888 20315 -10712
rect 15645 -15208 15785 -15032
rect 11115 -19528 11255 -19352
rect 6585 -23848 6725 -23672
rect 2055 -28168 2195 -27992
rect -2475 -32400 -2335 -32312
rect -165 -32400 -25 -32210
rect 2055 -32312 2075 -28168
rect 2175 -32312 2195 -28168
rect 4365 -28270 4505 -27890
rect 6585 -27992 6605 -23848
rect 6705 -27992 6725 -23848
rect 8895 -23950 9035 -23570
rect 11115 -23672 11135 -19528
rect 11235 -23672 11255 -19528
rect 13425 -19630 13565 -19250
rect 15645 -19352 15665 -15208
rect 15765 -19352 15785 -15208
rect 17955 -15310 18095 -14930
rect 20175 -15032 20195 -10888
rect 20295 -15032 20315 -10888
rect 22485 -10990 22625 -10610
rect 24705 -10712 24725 -6568
rect 24825 -10712 24845 -6568
rect 24705 -10888 24845 -10712
rect 20175 -15208 20315 -15032
rect 15645 -19528 15785 -19352
rect 11115 -23848 11255 -23672
rect 6585 -28168 6725 -27992
rect 2055 -32400 2195 -32312
rect 4365 -32400 4505 -32210
rect 6585 -32312 6605 -28168
rect 6705 -32312 6725 -28168
rect 8895 -28270 9035 -27890
rect 11115 -27992 11135 -23848
rect 11235 -27992 11255 -23848
rect 13425 -23950 13565 -23570
rect 15645 -23672 15665 -19528
rect 15765 -23672 15785 -19528
rect 17955 -19630 18095 -19250
rect 20175 -19352 20195 -15208
rect 20295 -19352 20315 -15208
rect 22485 -15310 22625 -14930
rect 24705 -15032 24725 -10888
rect 24825 -15032 24845 -10888
rect 24705 -15208 24845 -15032
rect 20175 -19528 20315 -19352
rect 15645 -23848 15785 -23672
rect 11115 -28168 11255 -27992
rect 6585 -32400 6725 -32312
rect 8895 -32400 9035 -32210
rect 11115 -32312 11135 -28168
rect 11235 -32312 11255 -28168
rect 13425 -28270 13565 -27890
rect 15645 -27992 15665 -23848
rect 15765 -27992 15785 -23848
rect 17955 -23950 18095 -23570
rect 20175 -23672 20195 -19528
rect 20295 -23672 20315 -19528
rect 22485 -19630 22625 -19250
rect 24705 -19352 24725 -15208
rect 24825 -19352 24845 -15208
rect 24705 -19528 24845 -19352
rect 20175 -23848 20315 -23672
rect 15645 -28168 15785 -27992
rect 11115 -32400 11255 -32312
rect 13425 -32400 13565 -32210
rect 15645 -32312 15665 -28168
rect 15765 -32312 15785 -28168
rect 17955 -28270 18095 -27890
rect 20175 -27992 20195 -23848
rect 20295 -27992 20315 -23848
rect 22485 -23950 22625 -23570
rect 24705 -23672 24725 -19528
rect 24825 -23672 24845 -19528
rect 24705 -23848 24845 -23672
rect 20175 -28168 20315 -27992
rect 15645 -32400 15785 -32312
rect 17955 -32400 18095 -32210
rect 20175 -32312 20195 -28168
rect 20295 -32312 20315 -28168
rect 22485 -28270 22625 -27890
rect 24705 -27992 24725 -23848
rect 24825 -27992 24845 -23848
rect 24705 -28168 24845 -27992
rect 20175 -32400 20315 -32312
rect 22485 -32400 22625 -32210
rect 24705 -32312 24725 -28168
rect 24825 -32312 24845 -28168
rect 24705 -32400 24845 -32312
<< properties >>
string parameters w 20.00 l 20.00 val 413.6 carea 1.00 cperi 0.17 nx 11 ny 15 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
