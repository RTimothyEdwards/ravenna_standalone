magic
tech EFXH018D
timestamp 1565723183
<< mimcap >>
rect -2180 42025 -180 42040
rect -2180 40055 -2165 42025
rect -195 40055 -180 42025
rect -2180 40040 -180 40055
rect 85 42025 2085 42040
rect 85 40055 100 42025
rect 2070 40055 2085 42025
rect 85 40040 2085 40055
rect -2180 39865 -180 39880
rect -2180 37895 -2165 39865
rect -195 37895 -180 39865
rect -2180 37880 -180 37895
rect 85 39865 2085 39880
rect 85 37895 100 39865
rect 2070 37895 2085 39865
rect 85 37880 2085 37895
rect -2180 37705 -180 37720
rect -2180 35735 -2165 37705
rect -195 35735 -180 37705
rect -2180 35720 -180 35735
rect 85 37705 2085 37720
rect 85 35735 100 37705
rect 2070 35735 2085 37705
rect 85 35720 2085 35735
rect -2180 35545 -180 35560
rect -2180 33575 -2165 35545
rect -195 33575 -180 35545
rect -2180 33560 -180 33575
rect 85 35545 2085 35560
rect 85 33575 100 35545
rect 2070 33575 2085 35545
rect 85 33560 2085 33575
rect -2180 33385 -180 33400
rect -2180 31415 -2165 33385
rect -195 31415 -180 33385
rect -2180 31400 -180 31415
rect 85 33385 2085 33400
rect 85 31415 100 33385
rect 2070 31415 2085 33385
rect 85 31400 2085 31415
rect -2180 31225 -180 31240
rect -2180 29255 -2165 31225
rect -195 29255 -180 31225
rect -2180 29240 -180 29255
rect 85 31225 2085 31240
rect 85 29255 100 31225
rect 2070 29255 2085 31225
rect 85 29240 2085 29255
rect -2180 29065 -180 29080
rect -2180 27095 -2165 29065
rect -195 27095 -180 29065
rect -2180 27080 -180 27095
rect 85 29065 2085 29080
rect 85 27095 100 29065
rect 2070 27095 2085 29065
rect 85 27080 2085 27095
rect -2180 26905 -180 26920
rect -2180 24935 -2165 26905
rect -195 24935 -180 26905
rect -2180 24920 -180 24935
rect 85 26905 2085 26920
rect 85 24935 100 26905
rect 2070 24935 2085 26905
rect 85 24920 2085 24935
rect -2180 24745 -180 24760
rect -2180 22775 -2165 24745
rect -195 22775 -180 24745
rect -2180 22760 -180 22775
rect 85 24745 2085 24760
rect 85 22775 100 24745
rect 2070 22775 2085 24745
rect 85 22760 2085 22775
rect -2180 22585 -180 22600
rect -2180 20615 -2165 22585
rect -195 20615 -180 22585
rect -2180 20600 -180 20615
rect 85 22585 2085 22600
rect 85 20615 100 22585
rect 2070 20615 2085 22585
rect 85 20600 2085 20615
rect -2180 20425 -180 20440
rect -2180 18455 -2165 20425
rect -195 18455 -180 20425
rect -2180 18440 -180 18455
rect 85 20425 2085 20440
rect 85 18455 100 20425
rect 2070 18455 2085 20425
rect 85 18440 2085 18455
rect -2180 18265 -180 18280
rect -2180 16295 -2165 18265
rect -195 16295 -180 18265
rect -2180 16280 -180 16295
rect 85 18265 2085 18280
rect 85 16295 100 18265
rect 2070 16295 2085 18265
rect 85 16280 2085 16295
rect -2180 16105 -180 16120
rect -2180 14135 -2165 16105
rect -195 14135 -180 16105
rect -2180 14120 -180 14135
rect 85 16105 2085 16120
rect 85 14135 100 16105
rect 2070 14135 2085 16105
rect 85 14120 2085 14135
rect -2180 13945 -180 13960
rect -2180 11975 -2165 13945
rect -195 11975 -180 13945
rect -2180 11960 -180 11975
rect 85 13945 2085 13960
rect 85 11975 100 13945
rect 2070 11975 2085 13945
rect 85 11960 2085 11975
rect -2180 11785 -180 11800
rect -2180 9815 -2165 11785
rect -195 9815 -180 11785
rect -2180 9800 -180 9815
rect 85 11785 2085 11800
rect 85 9815 100 11785
rect 2070 9815 2085 11785
rect 85 9800 2085 9815
rect -2180 9625 -180 9640
rect -2180 7655 -2165 9625
rect -195 7655 -180 9625
rect -2180 7640 -180 7655
rect 85 9625 2085 9640
rect 85 7655 100 9625
rect 2070 7655 2085 9625
rect 85 7640 2085 7655
rect -2180 7465 -180 7480
rect -2180 5495 -2165 7465
rect -195 5495 -180 7465
rect -2180 5480 -180 5495
rect 85 7465 2085 7480
rect 85 5495 100 7465
rect 2070 5495 2085 7465
rect 85 5480 2085 5495
rect -2180 5305 -180 5320
rect -2180 3335 -2165 5305
rect -195 3335 -180 5305
rect -2180 3320 -180 3335
rect 85 5305 2085 5320
rect 85 3335 100 5305
rect 2070 3335 2085 5305
rect 85 3320 2085 3335
rect -2180 3145 -180 3160
rect -2180 1175 -2165 3145
rect -195 1175 -180 3145
rect -2180 1160 -180 1175
rect 85 3145 2085 3160
rect 85 1175 100 3145
rect 2070 1175 2085 3145
rect 85 1160 2085 1175
rect -2180 985 -180 1000
rect -2180 -985 -2165 985
rect -195 -985 -180 985
rect -2180 -1000 -180 -985
rect 85 985 2085 1000
rect 85 -985 100 985
rect 2070 -985 2085 985
rect 85 -1000 2085 -985
rect -2180 -1175 -180 -1160
rect -2180 -3145 -2165 -1175
rect -195 -3145 -180 -1175
rect -2180 -3160 -180 -3145
rect 85 -1175 2085 -1160
rect 85 -3145 100 -1175
rect 2070 -3145 2085 -1175
rect 85 -3160 2085 -3145
rect -2180 -3335 -180 -3320
rect -2180 -5305 -2165 -3335
rect -195 -5305 -180 -3335
rect -2180 -5320 -180 -5305
rect 85 -3335 2085 -3320
rect 85 -5305 100 -3335
rect 2070 -5305 2085 -3335
rect 85 -5320 2085 -5305
rect -2180 -5495 -180 -5480
rect -2180 -7465 -2165 -5495
rect -195 -7465 -180 -5495
rect -2180 -7480 -180 -7465
rect 85 -5495 2085 -5480
rect 85 -7465 100 -5495
rect 2070 -7465 2085 -5495
rect 85 -7480 2085 -7465
rect -2180 -7655 -180 -7640
rect -2180 -9625 -2165 -7655
rect -195 -9625 -180 -7655
rect -2180 -9640 -180 -9625
rect 85 -7655 2085 -7640
rect 85 -9625 100 -7655
rect 2070 -9625 2085 -7655
rect 85 -9640 2085 -9625
rect -2180 -9815 -180 -9800
rect -2180 -11785 -2165 -9815
rect -195 -11785 -180 -9815
rect -2180 -11800 -180 -11785
rect 85 -9815 2085 -9800
rect 85 -11785 100 -9815
rect 2070 -11785 2085 -9815
rect 85 -11800 2085 -11785
rect -2180 -11975 -180 -11960
rect -2180 -13945 -2165 -11975
rect -195 -13945 -180 -11975
rect -2180 -13960 -180 -13945
rect 85 -11975 2085 -11960
rect 85 -13945 100 -11975
rect 2070 -13945 2085 -11975
rect 85 -13960 2085 -13945
rect -2180 -14135 -180 -14120
rect -2180 -16105 -2165 -14135
rect -195 -16105 -180 -14135
rect -2180 -16120 -180 -16105
rect 85 -14135 2085 -14120
rect 85 -16105 100 -14135
rect 2070 -16105 2085 -14135
rect 85 -16120 2085 -16105
rect -2180 -16295 -180 -16280
rect -2180 -18265 -2165 -16295
rect -195 -18265 -180 -16295
rect -2180 -18280 -180 -18265
rect 85 -16295 2085 -16280
rect 85 -18265 100 -16295
rect 2070 -18265 2085 -16295
rect 85 -18280 2085 -18265
rect -2180 -18455 -180 -18440
rect -2180 -20425 -2165 -18455
rect -195 -20425 -180 -18455
rect -2180 -20440 -180 -20425
rect 85 -18455 2085 -18440
rect 85 -20425 100 -18455
rect 2070 -20425 2085 -18455
rect 85 -20440 2085 -20425
rect -2180 -20615 -180 -20600
rect -2180 -22585 -2165 -20615
rect -195 -22585 -180 -20615
rect -2180 -22600 -180 -22585
rect 85 -20615 2085 -20600
rect 85 -22585 100 -20615
rect 2070 -22585 2085 -20615
rect 85 -22600 2085 -22585
rect -2180 -22775 -180 -22760
rect -2180 -24745 -2165 -22775
rect -195 -24745 -180 -22775
rect -2180 -24760 -180 -24745
rect 85 -22775 2085 -22760
rect 85 -24745 100 -22775
rect 2070 -24745 2085 -22775
rect 85 -24760 2085 -24745
rect -2180 -24935 -180 -24920
rect -2180 -26905 -2165 -24935
rect -195 -26905 -180 -24935
rect -2180 -26920 -180 -26905
rect 85 -24935 2085 -24920
rect 85 -26905 100 -24935
rect 2070 -26905 2085 -24935
rect 85 -26920 2085 -26905
rect -2180 -27095 -180 -27080
rect -2180 -29065 -2165 -27095
rect -195 -29065 -180 -27095
rect -2180 -29080 -180 -29065
rect 85 -27095 2085 -27080
rect 85 -29065 100 -27095
rect 2070 -29065 2085 -27095
rect 85 -29080 2085 -29065
rect -2180 -29255 -180 -29240
rect -2180 -31225 -2165 -29255
rect -195 -31225 -180 -29255
rect -2180 -31240 -180 -31225
rect 85 -29255 2085 -29240
rect 85 -31225 100 -29255
rect 2070 -31225 2085 -29255
rect 85 -31240 2085 -31225
rect -2180 -31415 -180 -31400
rect -2180 -33385 -2165 -31415
rect -195 -33385 -180 -31415
rect -2180 -33400 -180 -33385
rect 85 -31415 2085 -31400
rect 85 -33385 100 -31415
rect 2070 -33385 2085 -31415
rect 85 -33400 2085 -33385
rect -2180 -33575 -180 -33560
rect -2180 -35545 -2165 -33575
rect -195 -35545 -180 -33575
rect -2180 -35560 -180 -35545
rect 85 -33575 2085 -33560
rect 85 -35545 100 -33575
rect 2070 -35545 2085 -33575
rect 85 -35560 2085 -35545
rect -2180 -35735 -180 -35720
rect -2180 -37705 -2165 -35735
rect -195 -37705 -180 -35735
rect -2180 -37720 -180 -37705
rect 85 -35735 2085 -35720
rect 85 -37705 100 -35735
rect 2070 -37705 2085 -35735
rect 85 -37720 2085 -37705
rect -2180 -37895 -180 -37880
rect -2180 -39865 -2165 -37895
rect -195 -39865 -180 -37895
rect -2180 -39880 -180 -39865
rect 85 -37895 2085 -37880
rect 85 -39865 100 -37895
rect 2070 -39865 2085 -37895
rect 85 -39880 2085 -39865
rect -2180 -40055 -180 -40040
rect -2180 -42025 -2165 -40055
rect -195 -42025 -180 -40055
rect -2180 -42040 -180 -42025
rect 85 -40055 2085 -40040
rect 85 -42025 100 -40055
rect 2070 -42025 2085 -40055
rect 85 -42040 2085 -42025
<< mimcapcontact >>
rect -2165 40055 -195 42025
rect 100 40055 2070 42025
rect -2165 37895 -195 39865
rect 100 37895 2070 39865
rect -2165 35735 -195 37705
rect 100 35735 2070 37705
rect -2165 33575 -195 35545
rect 100 33575 2070 35545
rect -2165 31415 -195 33385
rect 100 31415 2070 33385
rect -2165 29255 -195 31225
rect 100 29255 2070 31225
rect -2165 27095 -195 29065
rect 100 27095 2070 29065
rect -2165 24935 -195 26905
rect 100 24935 2070 26905
rect -2165 22775 -195 24745
rect 100 22775 2070 24745
rect -2165 20615 -195 22585
rect 100 20615 2070 22585
rect -2165 18455 -195 20425
rect 100 18455 2070 20425
rect -2165 16295 -195 18265
rect 100 16295 2070 18265
rect -2165 14135 -195 16105
rect 100 14135 2070 16105
rect -2165 11975 -195 13945
rect 100 11975 2070 13945
rect -2165 9815 -195 11785
rect 100 9815 2070 11785
rect -2165 7655 -195 9625
rect 100 7655 2070 9625
rect -2165 5495 -195 7465
rect 100 5495 2070 7465
rect -2165 3335 -195 5305
rect 100 3335 2070 5305
rect -2165 1175 -195 3145
rect 100 1175 2070 3145
rect -2165 -985 -195 985
rect 100 -985 2070 985
rect -2165 -3145 -195 -1175
rect 100 -3145 2070 -1175
rect -2165 -5305 -195 -3335
rect 100 -5305 2070 -3335
rect -2165 -7465 -195 -5495
rect 100 -7465 2070 -5495
rect -2165 -9625 -195 -7655
rect 100 -9625 2070 -7655
rect -2165 -11785 -195 -9815
rect 100 -11785 2070 -9815
rect -2165 -13945 -195 -11975
rect 100 -13945 2070 -11975
rect -2165 -16105 -195 -14135
rect 100 -16105 2070 -14135
rect -2165 -18265 -195 -16295
rect 100 -18265 2070 -16295
rect -2165 -20425 -195 -18455
rect 100 -20425 2070 -18455
rect -2165 -22585 -195 -20615
rect 100 -22585 2070 -20615
rect -2165 -24745 -195 -22775
rect 100 -24745 2070 -22775
rect -2165 -26905 -195 -24935
rect 100 -26905 2070 -24935
rect -2165 -29065 -195 -27095
rect 100 -29065 2070 -27095
rect -2165 -31225 -195 -29255
rect 100 -31225 2070 -29255
rect -2165 -33385 -195 -31415
rect 100 -33385 2070 -31415
rect -2165 -35545 -195 -33575
rect 100 -35545 2070 -33575
rect -2165 -37705 -195 -35735
rect 100 -37705 2070 -35735
rect -2165 -39865 -195 -37895
rect 100 -39865 2070 -37895
rect -2165 -42025 -195 -40055
rect 100 -42025 2070 -40055
<< metal4 >>
rect -2230 42076 -35 42090
rect -2230 42040 -95 42076
rect -2230 40040 -2180 42040
rect -180 40040 -95 42040
rect -2230 40004 -95 40040
rect -45 40004 -35 42076
rect -2230 39990 -35 40004
rect 35 42076 2230 42090
rect 35 42040 2170 42076
rect 35 40040 85 42040
rect 2085 40040 2170 42040
rect 35 40004 2170 40040
rect 2220 40004 2230 42076
rect 35 39990 2230 40004
rect -2230 39916 -35 39930
rect -2230 39880 -95 39916
rect -2230 37880 -2180 39880
rect -180 37880 -95 39880
rect -2230 37844 -95 37880
rect -45 37844 -35 39916
rect -2230 37830 -35 37844
rect 35 39916 2230 39930
rect 35 39880 2170 39916
rect 35 37880 85 39880
rect 2085 37880 2170 39880
rect 35 37844 2170 37880
rect 2220 37844 2230 39916
rect 35 37830 2230 37844
rect -2230 37756 -35 37770
rect -2230 37720 -95 37756
rect -2230 35720 -2180 37720
rect -180 35720 -95 37720
rect -2230 35684 -95 35720
rect -45 35684 -35 37756
rect -2230 35670 -35 35684
rect 35 37756 2230 37770
rect 35 37720 2170 37756
rect 35 35720 85 37720
rect 2085 35720 2170 37720
rect 35 35684 2170 35720
rect 2220 35684 2230 37756
rect 35 35670 2230 35684
rect -2230 35596 -35 35610
rect -2230 35560 -95 35596
rect -2230 33560 -2180 35560
rect -180 33560 -95 35560
rect -2230 33524 -95 33560
rect -45 33524 -35 35596
rect -2230 33510 -35 33524
rect 35 35596 2230 35610
rect 35 35560 2170 35596
rect 35 33560 85 35560
rect 2085 33560 2170 35560
rect 35 33524 2170 33560
rect 2220 33524 2230 35596
rect 35 33510 2230 33524
rect -2230 33436 -35 33450
rect -2230 33400 -95 33436
rect -2230 31400 -2180 33400
rect -180 31400 -95 33400
rect -2230 31364 -95 31400
rect -45 31364 -35 33436
rect -2230 31350 -35 31364
rect 35 33436 2230 33450
rect 35 33400 2170 33436
rect 35 31400 85 33400
rect 2085 31400 2170 33400
rect 35 31364 2170 31400
rect 2220 31364 2230 33436
rect 35 31350 2230 31364
rect -2230 31276 -35 31290
rect -2230 31240 -95 31276
rect -2230 29240 -2180 31240
rect -180 29240 -95 31240
rect -2230 29204 -95 29240
rect -45 29204 -35 31276
rect -2230 29190 -35 29204
rect 35 31276 2230 31290
rect 35 31240 2170 31276
rect 35 29240 85 31240
rect 2085 29240 2170 31240
rect 35 29204 2170 29240
rect 2220 29204 2230 31276
rect 35 29190 2230 29204
rect -2230 29116 -35 29130
rect -2230 29080 -95 29116
rect -2230 27080 -2180 29080
rect -180 27080 -95 29080
rect -2230 27044 -95 27080
rect -45 27044 -35 29116
rect -2230 27030 -35 27044
rect 35 29116 2230 29130
rect 35 29080 2170 29116
rect 35 27080 85 29080
rect 2085 27080 2170 29080
rect 35 27044 2170 27080
rect 2220 27044 2230 29116
rect 35 27030 2230 27044
rect -2230 26956 -35 26970
rect -2230 26920 -95 26956
rect -2230 24920 -2180 26920
rect -180 24920 -95 26920
rect -2230 24884 -95 24920
rect -45 24884 -35 26956
rect -2230 24870 -35 24884
rect 35 26956 2230 26970
rect 35 26920 2170 26956
rect 35 24920 85 26920
rect 2085 24920 2170 26920
rect 35 24884 2170 24920
rect 2220 24884 2230 26956
rect 35 24870 2230 24884
rect -2230 24796 -35 24810
rect -2230 24760 -95 24796
rect -2230 22760 -2180 24760
rect -180 22760 -95 24760
rect -2230 22724 -95 22760
rect -45 22724 -35 24796
rect -2230 22710 -35 22724
rect 35 24796 2230 24810
rect 35 24760 2170 24796
rect 35 22760 85 24760
rect 2085 22760 2170 24760
rect 35 22724 2170 22760
rect 2220 22724 2230 24796
rect 35 22710 2230 22724
rect -2230 22636 -35 22650
rect -2230 22600 -95 22636
rect -2230 20600 -2180 22600
rect -180 20600 -95 22600
rect -2230 20564 -95 20600
rect -45 20564 -35 22636
rect -2230 20550 -35 20564
rect 35 22636 2230 22650
rect 35 22600 2170 22636
rect 35 20600 85 22600
rect 2085 20600 2170 22600
rect 35 20564 2170 20600
rect 2220 20564 2230 22636
rect 35 20550 2230 20564
rect -2230 20476 -35 20490
rect -2230 20440 -95 20476
rect -2230 18440 -2180 20440
rect -180 18440 -95 20440
rect -2230 18404 -95 18440
rect -45 18404 -35 20476
rect -2230 18390 -35 18404
rect 35 20476 2230 20490
rect 35 20440 2170 20476
rect 35 18440 85 20440
rect 2085 18440 2170 20440
rect 35 18404 2170 18440
rect 2220 18404 2230 20476
rect 35 18390 2230 18404
rect -2230 18316 -35 18330
rect -2230 18280 -95 18316
rect -2230 16280 -2180 18280
rect -180 16280 -95 18280
rect -2230 16244 -95 16280
rect -45 16244 -35 18316
rect -2230 16230 -35 16244
rect 35 18316 2230 18330
rect 35 18280 2170 18316
rect 35 16280 85 18280
rect 2085 16280 2170 18280
rect 35 16244 2170 16280
rect 2220 16244 2230 18316
rect 35 16230 2230 16244
rect -2230 16156 -35 16170
rect -2230 16120 -95 16156
rect -2230 14120 -2180 16120
rect -180 14120 -95 16120
rect -2230 14084 -95 14120
rect -45 14084 -35 16156
rect -2230 14070 -35 14084
rect 35 16156 2230 16170
rect 35 16120 2170 16156
rect 35 14120 85 16120
rect 2085 14120 2170 16120
rect 35 14084 2170 14120
rect 2220 14084 2230 16156
rect 35 14070 2230 14084
rect -2230 13996 -35 14010
rect -2230 13960 -95 13996
rect -2230 11960 -2180 13960
rect -180 11960 -95 13960
rect -2230 11924 -95 11960
rect -45 11924 -35 13996
rect -2230 11910 -35 11924
rect 35 13996 2230 14010
rect 35 13960 2170 13996
rect 35 11960 85 13960
rect 2085 11960 2170 13960
rect 35 11924 2170 11960
rect 2220 11924 2230 13996
rect 35 11910 2230 11924
rect -2230 11836 -35 11850
rect -2230 11800 -95 11836
rect -2230 9800 -2180 11800
rect -180 9800 -95 11800
rect -2230 9764 -95 9800
rect -45 9764 -35 11836
rect -2230 9750 -35 9764
rect 35 11836 2230 11850
rect 35 11800 2170 11836
rect 35 9800 85 11800
rect 2085 9800 2170 11800
rect 35 9764 2170 9800
rect 2220 9764 2230 11836
rect 35 9750 2230 9764
rect -2230 9676 -35 9690
rect -2230 9640 -95 9676
rect -2230 7640 -2180 9640
rect -180 7640 -95 9640
rect -2230 7604 -95 7640
rect -45 7604 -35 9676
rect -2230 7590 -35 7604
rect 35 9676 2230 9690
rect 35 9640 2170 9676
rect 35 7640 85 9640
rect 2085 7640 2170 9640
rect 35 7604 2170 7640
rect 2220 7604 2230 9676
rect 35 7590 2230 7604
rect -2230 7516 -35 7530
rect -2230 7480 -95 7516
rect -2230 5480 -2180 7480
rect -180 5480 -95 7480
rect -2230 5444 -95 5480
rect -45 5444 -35 7516
rect -2230 5430 -35 5444
rect 35 7516 2230 7530
rect 35 7480 2170 7516
rect 35 5480 85 7480
rect 2085 5480 2170 7480
rect 35 5444 2170 5480
rect 2220 5444 2230 7516
rect 35 5430 2230 5444
rect -2230 5356 -35 5370
rect -2230 5320 -95 5356
rect -2230 3320 -2180 5320
rect -180 3320 -95 5320
rect -2230 3284 -95 3320
rect -45 3284 -35 5356
rect -2230 3270 -35 3284
rect 35 5356 2230 5370
rect 35 5320 2170 5356
rect 35 3320 85 5320
rect 2085 3320 2170 5320
rect 35 3284 2170 3320
rect 2220 3284 2230 5356
rect 35 3270 2230 3284
rect -2230 3196 -35 3210
rect -2230 3160 -95 3196
rect -2230 1160 -2180 3160
rect -180 1160 -95 3160
rect -2230 1124 -95 1160
rect -45 1124 -35 3196
rect -2230 1110 -35 1124
rect 35 3196 2230 3210
rect 35 3160 2170 3196
rect 35 1160 85 3160
rect 2085 1160 2170 3160
rect 35 1124 2170 1160
rect 2220 1124 2230 3196
rect 35 1110 2230 1124
rect -2230 1036 -35 1050
rect -2230 1000 -95 1036
rect -2230 -1000 -2180 1000
rect -180 -1000 -95 1000
rect -2230 -1036 -95 -1000
rect -45 -1036 -35 1036
rect -2230 -1050 -35 -1036
rect 35 1036 2230 1050
rect 35 1000 2170 1036
rect 35 -1000 85 1000
rect 2085 -1000 2170 1000
rect 35 -1036 2170 -1000
rect 2220 -1036 2230 1036
rect 35 -1050 2230 -1036
rect -2230 -1124 -35 -1110
rect -2230 -1160 -95 -1124
rect -2230 -3160 -2180 -1160
rect -180 -3160 -95 -1160
rect -2230 -3196 -95 -3160
rect -45 -3196 -35 -1124
rect -2230 -3210 -35 -3196
rect 35 -1124 2230 -1110
rect 35 -1160 2170 -1124
rect 35 -3160 85 -1160
rect 2085 -3160 2170 -1160
rect 35 -3196 2170 -3160
rect 2220 -3196 2230 -1124
rect 35 -3210 2230 -3196
rect -2230 -3284 -35 -3270
rect -2230 -3320 -95 -3284
rect -2230 -5320 -2180 -3320
rect -180 -5320 -95 -3320
rect -2230 -5356 -95 -5320
rect -45 -5356 -35 -3284
rect -2230 -5370 -35 -5356
rect 35 -3284 2230 -3270
rect 35 -3320 2170 -3284
rect 35 -5320 85 -3320
rect 2085 -5320 2170 -3320
rect 35 -5356 2170 -5320
rect 2220 -5356 2230 -3284
rect 35 -5370 2230 -5356
rect -2230 -5444 -35 -5430
rect -2230 -5480 -95 -5444
rect -2230 -7480 -2180 -5480
rect -180 -7480 -95 -5480
rect -2230 -7516 -95 -7480
rect -45 -7516 -35 -5444
rect -2230 -7530 -35 -7516
rect 35 -5444 2230 -5430
rect 35 -5480 2170 -5444
rect 35 -7480 85 -5480
rect 2085 -7480 2170 -5480
rect 35 -7516 2170 -7480
rect 2220 -7516 2230 -5444
rect 35 -7530 2230 -7516
rect -2230 -7604 -35 -7590
rect -2230 -7640 -95 -7604
rect -2230 -9640 -2180 -7640
rect -180 -9640 -95 -7640
rect -2230 -9676 -95 -9640
rect -45 -9676 -35 -7604
rect -2230 -9690 -35 -9676
rect 35 -7604 2230 -7590
rect 35 -7640 2170 -7604
rect 35 -9640 85 -7640
rect 2085 -9640 2170 -7640
rect 35 -9676 2170 -9640
rect 2220 -9676 2230 -7604
rect 35 -9690 2230 -9676
rect -2230 -9764 -35 -9750
rect -2230 -9800 -95 -9764
rect -2230 -11800 -2180 -9800
rect -180 -11800 -95 -9800
rect -2230 -11836 -95 -11800
rect -45 -11836 -35 -9764
rect -2230 -11850 -35 -11836
rect 35 -9764 2230 -9750
rect 35 -9800 2170 -9764
rect 35 -11800 85 -9800
rect 2085 -11800 2170 -9800
rect 35 -11836 2170 -11800
rect 2220 -11836 2230 -9764
rect 35 -11850 2230 -11836
rect -2230 -11924 -35 -11910
rect -2230 -11960 -95 -11924
rect -2230 -13960 -2180 -11960
rect -180 -13960 -95 -11960
rect -2230 -13996 -95 -13960
rect -45 -13996 -35 -11924
rect -2230 -14010 -35 -13996
rect 35 -11924 2230 -11910
rect 35 -11960 2170 -11924
rect 35 -13960 85 -11960
rect 2085 -13960 2170 -11960
rect 35 -13996 2170 -13960
rect 2220 -13996 2230 -11924
rect 35 -14010 2230 -13996
rect -2230 -14084 -35 -14070
rect -2230 -14120 -95 -14084
rect -2230 -16120 -2180 -14120
rect -180 -16120 -95 -14120
rect -2230 -16156 -95 -16120
rect -45 -16156 -35 -14084
rect -2230 -16170 -35 -16156
rect 35 -14084 2230 -14070
rect 35 -14120 2170 -14084
rect 35 -16120 85 -14120
rect 2085 -16120 2170 -14120
rect 35 -16156 2170 -16120
rect 2220 -16156 2230 -14084
rect 35 -16170 2230 -16156
rect -2230 -16244 -35 -16230
rect -2230 -16280 -95 -16244
rect -2230 -18280 -2180 -16280
rect -180 -18280 -95 -16280
rect -2230 -18316 -95 -18280
rect -45 -18316 -35 -16244
rect -2230 -18330 -35 -18316
rect 35 -16244 2230 -16230
rect 35 -16280 2170 -16244
rect 35 -18280 85 -16280
rect 2085 -18280 2170 -16280
rect 35 -18316 2170 -18280
rect 2220 -18316 2230 -16244
rect 35 -18330 2230 -18316
rect -2230 -18404 -35 -18390
rect -2230 -18440 -95 -18404
rect -2230 -20440 -2180 -18440
rect -180 -20440 -95 -18440
rect -2230 -20476 -95 -20440
rect -45 -20476 -35 -18404
rect -2230 -20490 -35 -20476
rect 35 -18404 2230 -18390
rect 35 -18440 2170 -18404
rect 35 -20440 85 -18440
rect 2085 -20440 2170 -18440
rect 35 -20476 2170 -20440
rect 2220 -20476 2230 -18404
rect 35 -20490 2230 -20476
rect -2230 -20564 -35 -20550
rect -2230 -20600 -95 -20564
rect -2230 -22600 -2180 -20600
rect -180 -22600 -95 -20600
rect -2230 -22636 -95 -22600
rect -45 -22636 -35 -20564
rect -2230 -22650 -35 -22636
rect 35 -20564 2230 -20550
rect 35 -20600 2170 -20564
rect 35 -22600 85 -20600
rect 2085 -22600 2170 -20600
rect 35 -22636 2170 -22600
rect 2220 -22636 2230 -20564
rect 35 -22650 2230 -22636
rect -2230 -22724 -35 -22710
rect -2230 -22760 -95 -22724
rect -2230 -24760 -2180 -22760
rect -180 -24760 -95 -22760
rect -2230 -24796 -95 -24760
rect -45 -24796 -35 -22724
rect -2230 -24810 -35 -24796
rect 35 -22724 2230 -22710
rect 35 -22760 2170 -22724
rect 35 -24760 85 -22760
rect 2085 -24760 2170 -22760
rect 35 -24796 2170 -24760
rect 2220 -24796 2230 -22724
rect 35 -24810 2230 -24796
rect -2230 -24884 -35 -24870
rect -2230 -24920 -95 -24884
rect -2230 -26920 -2180 -24920
rect -180 -26920 -95 -24920
rect -2230 -26956 -95 -26920
rect -45 -26956 -35 -24884
rect -2230 -26970 -35 -26956
rect 35 -24884 2230 -24870
rect 35 -24920 2170 -24884
rect 35 -26920 85 -24920
rect 2085 -26920 2170 -24920
rect 35 -26956 2170 -26920
rect 2220 -26956 2230 -24884
rect 35 -26970 2230 -26956
rect -2230 -27044 -35 -27030
rect -2230 -27080 -95 -27044
rect -2230 -29080 -2180 -27080
rect -180 -29080 -95 -27080
rect -2230 -29116 -95 -29080
rect -45 -29116 -35 -27044
rect -2230 -29130 -35 -29116
rect 35 -27044 2230 -27030
rect 35 -27080 2170 -27044
rect 35 -29080 85 -27080
rect 2085 -29080 2170 -27080
rect 35 -29116 2170 -29080
rect 2220 -29116 2230 -27044
rect 35 -29130 2230 -29116
rect -2230 -29204 -35 -29190
rect -2230 -29240 -95 -29204
rect -2230 -31240 -2180 -29240
rect -180 -31240 -95 -29240
rect -2230 -31276 -95 -31240
rect -45 -31276 -35 -29204
rect -2230 -31290 -35 -31276
rect 35 -29204 2230 -29190
rect 35 -29240 2170 -29204
rect 35 -31240 85 -29240
rect 2085 -31240 2170 -29240
rect 35 -31276 2170 -31240
rect 2220 -31276 2230 -29204
rect 35 -31290 2230 -31276
rect -2230 -31364 -35 -31350
rect -2230 -31400 -95 -31364
rect -2230 -33400 -2180 -31400
rect -180 -33400 -95 -31400
rect -2230 -33436 -95 -33400
rect -45 -33436 -35 -31364
rect -2230 -33450 -35 -33436
rect 35 -31364 2230 -31350
rect 35 -31400 2170 -31364
rect 35 -33400 85 -31400
rect 2085 -33400 2170 -31400
rect 35 -33436 2170 -33400
rect 2220 -33436 2230 -31364
rect 35 -33450 2230 -33436
rect -2230 -33524 -35 -33510
rect -2230 -33560 -95 -33524
rect -2230 -35560 -2180 -33560
rect -180 -35560 -95 -33560
rect -2230 -35596 -95 -35560
rect -45 -35596 -35 -33524
rect -2230 -35610 -35 -35596
rect 35 -33524 2230 -33510
rect 35 -33560 2170 -33524
rect 35 -35560 85 -33560
rect 2085 -35560 2170 -33560
rect 35 -35596 2170 -35560
rect 2220 -35596 2230 -33524
rect 35 -35610 2230 -35596
rect -2230 -35684 -35 -35670
rect -2230 -35720 -95 -35684
rect -2230 -37720 -2180 -35720
rect -180 -37720 -95 -35720
rect -2230 -37756 -95 -37720
rect -45 -37756 -35 -35684
rect -2230 -37770 -35 -37756
rect 35 -35684 2230 -35670
rect 35 -35720 2170 -35684
rect 35 -37720 85 -35720
rect 2085 -37720 2170 -35720
rect 35 -37756 2170 -37720
rect 2220 -37756 2230 -35684
rect 35 -37770 2230 -37756
rect -2230 -37844 -35 -37830
rect -2230 -37880 -95 -37844
rect -2230 -39880 -2180 -37880
rect -180 -39880 -95 -37880
rect -2230 -39916 -95 -39880
rect -45 -39916 -35 -37844
rect -2230 -39930 -35 -39916
rect 35 -37844 2230 -37830
rect 35 -37880 2170 -37844
rect 35 -39880 85 -37880
rect 2085 -39880 2170 -37880
rect 35 -39916 2170 -39880
rect 2220 -39916 2230 -37844
rect 35 -39930 2230 -39916
rect -2230 -40004 -35 -39990
rect -2230 -40040 -95 -40004
rect -2230 -42040 -2180 -40040
rect -180 -42040 -95 -40040
rect -2230 -42076 -95 -42040
rect -45 -42076 -35 -40004
rect -2230 -42090 -35 -42076
rect 35 -40004 2230 -39990
rect 35 -40040 2170 -40004
rect 35 -42040 85 -40040
rect 2085 -42040 2170 -40040
rect 35 -42076 2170 -42040
rect 2220 -42076 2230 -40004
rect 35 -42090 2230 -42076
<< viatp >>
rect -95 40004 -45 42076
rect 2170 40004 2220 42076
rect -95 37844 -45 39916
rect 2170 37844 2220 39916
rect -95 35684 -45 37756
rect 2170 35684 2220 37756
rect -95 33524 -45 35596
rect 2170 33524 2220 35596
rect -95 31364 -45 33436
rect 2170 31364 2220 33436
rect -95 29204 -45 31276
rect 2170 29204 2220 31276
rect -95 27044 -45 29116
rect 2170 27044 2220 29116
rect -95 24884 -45 26956
rect 2170 24884 2220 26956
rect -95 22724 -45 24796
rect 2170 22724 2220 24796
rect -95 20564 -45 22636
rect 2170 20564 2220 22636
rect -95 18404 -45 20476
rect 2170 18404 2220 20476
rect -95 16244 -45 18316
rect 2170 16244 2220 18316
rect -95 14084 -45 16156
rect 2170 14084 2220 16156
rect -95 11924 -45 13996
rect 2170 11924 2220 13996
rect -95 9764 -45 11836
rect 2170 9764 2220 11836
rect -95 7604 -45 9676
rect 2170 7604 2220 9676
rect -95 5444 -45 7516
rect 2170 5444 2220 7516
rect -95 3284 -45 5356
rect 2170 3284 2220 5356
rect -95 1124 -45 3196
rect 2170 1124 2220 3196
rect -95 -1036 -45 1036
rect 2170 -1036 2220 1036
rect -95 -3196 -45 -1124
rect 2170 -3196 2220 -1124
rect -95 -5356 -45 -3284
rect 2170 -5356 2220 -3284
rect -95 -7516 -45 -5444
rect 2170 -7516 2220 -5444
rect -95 -9676 -45 -7604
rect 2170 -9676 2220 -7604
rect -95 -11836 -45 -9764
rect 2170 -11836 2220 -9764
rect -95 -13996 -45 -11924
rect 2170 -13996 2220 -11924
rect -95 -16156 -45 -14084
rect 2170 -16156 2220 -14084
rect -95 -18316 -45 -16244
rect 2170 -18316 2220 -16244
rect -95 -20476 -45 -18404
rect 2170 -20476 2220 -18404
rect -95 -22636 -45 -20564
rect 2170 -22636 2220 -20564
rect -95 -24796 -45 -22724
rect 2170 -24796 2220 -22724
rect -95 -26956 -45 -24884
rect 2170 -26956 2220 -24884
rect -95 -29116 -45 -27044
rect 2170 -29116 2220 -27044
rect -95 -31276 -45 -29204
rect 2170 -31276 2220 -29204
rect -95 -33436 -45 -31364
rect 2170 -33436 2220 -31364
rect -95 -35596 -45 -33524
rect 2170 -35596 2220 -33524
rect -95 -37756 -45 -35684
rect 2170 -37756 2220 -35684
rect -95 -39916 -45 -37844
rect 2170 -39916 2220 -37844
rect -95 -42076 -45 -40004
rect 2170 -42076 2220 -40004
<< metaltp >>
rect -1215 42025 -1145 42120
rect -105 42076 -35 42120
rect -1215 39865 -1145 40055
rect -105 40004 -95 42076
rect -45 40004 -35 42076
rect 1050 42025 1120 42120
rect 2160 42076 2230 42120
rect -105 39916 -35 40004
rect -1215 37705 -1145 37895
rect -105 37844 -95 39916
rect -45 37844 -35 39916
rect 1050 39865 1120 40055
rect 2160 40004 2170 42076
rect 2220 40004 2230 42076
rect 2160 39916 2230 40004
rect -105 37756 -35 37844
rect -1215 35545 -1145 35735
rect -105 35684 -95 37756
rect -45 35684 -35 37756
rect 1050 37705 1120 37895
rect 2160 37844 2170 39916
rect 2220 37844 2230 39916
rect 2160 37756 2230 37844
rect -105 35596 -35 35684
rect -1215 33385 -1145 33575
rect -105 33524 -95 35596
rect -45 33524 -35 35596
rect 1050 35545 1120 35735
rect 2160 35684 2170 37756
rect 2220 35684 2230 37756
rect 2160 35596 2230 35684
rect -105 33436 -35 33524
rect -1215 31225 -1145 31415
rect -105 31364 -95 33436
rect -45 31364 -35 33436
rect 1050 33385 1120 33575
rect 2160 33524 2170 35596
rect 2220 33524 2230 35596
rect 2160 33436 2230 33524
rect -105 31276 -35 31364
rect -1215 29065 -1145 29255
rect -105 29204 -95 31276
rect -45 29204 -35 31276
rect 1050 31225 1120 31415
rect 2160 31364 2170 33436
rect 2220 31364 2230 33436
rect 2160 31276 2230 31364
rect -105 29116 -35 29204
rect -1215 26905 -1145 27095
rect -105 27044 -95 29116
rect -45 27044 -35 29116
rect 1050 29065 1120 29255
rect 2160 29204 2170 31276
rect 2220 29204 2230 31276
rect 2160 29116 2230 29204
rect -105 26956 -35 27044
rect -1215 24745 -1145 24935
rect -105 24884 -95 26956
rect -45 24884 -35 26956
rect 1050 26905 1120 27095
rect 2160 27044 2170 29116
rect 2220 27044 2230 29116
rect 2160 26956 2230 27044
rect -105 24796 -35 24884
rect -1215 22585 -1145 22775
rect -105 22724 -95 24796
rect -45 22724 -35 24796
rect 1050 24745 1120 24935
rect 2160 24884 2170 26956
rect 2220 24884 2230 26956
rect 2160 24796 2230 24884
rect -105 22636 -35 22724
rect -1215 20425 -1145 20615
rect -105 20564 -95 22636
rect -45 20564 -35 22636
rect 1050 22585 1120 22775
rect 2160 22724 2170 24796
rect 2220 22724 2230 24796
rect 2160 22636 2230 22724
rect -105 20476 -35 20564
rect -1215 18265 -1145 18455
rect -105 18404 -95 20476
rect -45 18404 -35 20476
rect 1050 20425 1120 20615
rect 2160 20564 2170 22636
rect 2220 20564 2230 22636
rect 2160 20476 2230 20564
rect -105 18316 -35 18404
rect -1215 16105 -1145 16295
rect -105 16244 -95 18316
rect -45 16244 -35 18316
rect 1050 18265 1120 18455
rect 2160 18404 2170 20476
rect 2220 18404 2230 20476
rect 2160 18316 2230 18404
rect -105 16156 -35 16244
rect -1215 13945 -1145 14135
rect -105 14084 -95 16156
rect -45 14084 -35 16156
rect 1050 16105 1120 16295
rect 2160 16244 2170 18316
rect 2220 16244 2230 18316
rect 2160 16156 2230 16244
rect -105 13996 -35 14084
rect -1215 11785 -1145 11975
rect -105 11924 -95 13996
rect -45 11924 -35 13996
rect 1050 13945 1120 14135
rect 2160 14084 2170 16156
rect 2220 14084 2230 16156
rect 2160 13996 2230 14084
rect -105 11836 -35 11924
rect -1215 9625 -1145 9815
rect -105 9764 -95 11836
rect -45 9764 -35 11836
rect 1050 11785 1120 11975
rect 2160 11924 2170 13996
rect 2220 11924 2230 13996
rect 2160 11836 2230 11924
rect -105 9676 -35 9764
rect -1215 7465 -1145 7655
rect -105 7604 -95 9676
rect -45 7604 -35 9676
rect 1050 9625 1120 9815
rect 2160 9764 2170 11836
rect 2220 9764 2230 11836
rect 2160 9676 2230 9764
rect -105 7516 -35 7604
rect -1215 5305 -1145 5495
rect -105 5444 -95 7516
rect -45 5444 -35 7516
rect 1050 7465 1120 7655
rect 2160 7604 2170 9676
rect 2220 7604 2230 9676
rect 2160 7516 2230 7604
rect -105 5356 -35 5444
rect -1215 3145 -1145 3335
rect -105 3284 -95 5356
rect -45 3284 -35 5356
rect 1050 5305 1120 5495
rect 2160 5444 2170 7516
rect 2220 5444 2230 7516
rect 2160 5356 2230 5444
rect -105 3196 -35 3284
rect -1215 985 -1145 1175
rect -105 1124 -95 3196
rect -45 1124 -35 3196
rect 1050 3145 1120 3335
rect 2160 3284 2170 5356
rect 2220 3284 2230 5356
rect 2160 3196 2230 3284
rect -105 1036 -35 1124
rect -1215 -1175 -1145 -985
rect -105 -1036 -95 1036
rect -45 -1036 -35 1036
rect 1050 985 1120 1175
rect 2160 1124 2170 3196
rect 2220 1124 2230 3196
rect 2160 1036 2230 1124
rect -105 -1124 -35 -1036
rect -1215 -3335 -1145 -3145
rect -105 -3196 -95 -1124
rect -45 -3196 -35 -1124
rect 1050 -1175 1120 -985
rect 2160 -1036 2170 1036
rect 2220 -1036 2230 1036
rect 2160 -1124 2230 -1036
rect -105 -3284 -35 -3196
rect -1215 -5495 -1145 -5305
rect -105 -5356 -95 -3284
rect -45 -5356 -35 -3284
rect 1050 -3335 1120 -3145
rect 2160 -3196 2170 -1124
rect 2220 -3196 2230 -1124
rect 2160 -3284 2230 -3196
rect -105 -5444 -35 -5356
rect -1215 -7655 -1145 -7465
rect -105 -7516 -95 -5444
rect -45 -7516 -35 -5444
rect 1050 -5495 1120 -5305
rect 2160 -5356 2170 -3284
rect 2220 -5356 2230 -3284
rect 2160 -5444 2230 -5356
rect -105 -7604 -35 -7516
rect -1215 -9815 -1145 -9625
rect -105 -9676 -95 -7604
rect -45 -9676 -35 -7604
rect 1050 -7655 1120 -7465
rect 2160 -7516 2170 -5444
rect 2220 -7516 2230 -5444
rect 2160 -7604 2230 -7516
rect -105 -9764 -35 -9676
rect -1215 -11975 -1145 -11785
rect -105 -11836 -95 -9764
rect -45 -11836 -35 -9764
rect 1050 -9815 1120 -9625
rect 2160 -9676 2170 -7604
rect 2220 -9676 2230 -7604
rect 2160 -9764 2230 -9676
rect -105 -11924 -35 -11836
rect -1215 -14135 -1145 -13945
rect -105 -13996 -95 -11924
rect -45 -13996 -35 -11924
rect 1050 -11975 1120 -11785
rect 2160 -11836 2170 -9764
rect 2220 -11836 2230 -9764
rect 2160 -11924 2230 -11836
rect -105 -14084 -35 -13996
rect -1215 -16295 -1145 -16105
rect -105 -16156 -95 -14084
rect -45 -16156 -35 -14084
rect 1050 -14135 1120 -13945
rect 2160 -13996 2170 -11924
rect 2220 -13996 2230 -11924
rect 2160 -14084 2230 -13996
rect -105 -16244 -35 -16156
rect -1215 -18455 -1145 -18265
rect -105 -18316 -95 -16244
rect -45 -18316 -35 -16244
rect 1050 -16295 1120 -16105
rect 2160 -16156 2170 -14084
rect 2220 -16156 2230 -14084
rect 2160 -16244 2230 -16156
rect -105 -18404 -35 -18316
rect -1215 -20615 -1145 -20425
rect -105 -20476 -95 -18404
rect -45 -20476 -35 -18404
rect 1050 -18455 1120 -18265
rect 2160 -18316 2170 -16244
rect 2220 -18316 2230 -16244
rect 2160 -18404 2230 -18316
rect -105 -20564 -35 -20476
rect -1215 -22775 -1145 -22585
rect -105 -22636 -95 -20564
rect -45 -22636 -35 -20564
rect 1050 -20615 1120 -20425
rect 2160 -20476 2170 -18404
rect 2220 -20476 2230 -18404
rect 2160 -20564 2230 -20476
rect -105 -22724 -35 -22636
rect -1215 -24935 -1145 -24745
rect -105 -24796 -95 -22724
rect -45 -24796 -35 -22724
rect 1050 -22775 1120 -22585
rect 2160 -22636 2170 -20564
rect 2220 -22636 2230 -20564
rect 2160 -22724 2230 -22636
rect -105 -24884 -35 -24796
rect -1215 -27095 -1145 -26905
rect -105 -26956 -95 -24884
rect -45 -26956 -35 -24884
rect 1050 -24935 1120 -24745
rect 2160 -24796 2170 -22724
rect 2220 -24796 2230 -22724
rect 2160 -24884 2230 -24796
rect -105 -27044 -35 -26956
rect -1215 -29255 -1145 -29065
rect -105 -29116 -95 -27044
rect -45 -29116 -35 -27044
rect 1050 -27095 1120 -26905
rect 2160 -26956 2170 -24884
rect 2220 -26956 2230 -24884
rect 2160 -27044 2230 -26956
rect -105 -29204 -35 -29116
rect -1215 -31415 -1145 -31225
rect -105 -31276 -95 -29204
rect -45 -31276 -35 -29204
rect 1050 -29255 1120 -29065
rect 2160 -29116 2170 -27044
rect 2220 -29116 2230 -27044
rect 2160 -29204 2230 -29116
rect -105 -31364 -35 -31276
rect -1215 -33575 -1145 -33385
rect -105 -33436 -95 -31364
rect -45 -33436 -35 -31364
rect 1050 -31415 1120 -31225
rect 2160 -31276 2170 -29204
rect 2220 -31276 2230 -29204
rect 2160 -31364 2230 -31276
rect -105 -33524 -35 -33436
rect -1215 -35735 -1145 -35545
rect -105 -35596 -95 -33524
rect -45 -35596 -35 -33524
rect 1050 -33575 1120 -33385
rect 2160 -33436 2170 -31364
rect 2220 -33436 2230 -31364
rect 2160 -33524 2230 -33436
rect -105 -35684 -35 -35596
rect -1215 -37895 -1145 -37705
rect -105 -37756 -95 -35684
rect -45 -37756 -35 -35684
rect 1050 -35735 1120 -35545
rect 2160 -35596 2170 -33524
rect 2220 -35596 2230 -33524
rect 2160 -35684 2230 -35596
rect -105 -37844 -35 -37756
rect -1215 -40055 -1145 -39865
rect -105 -39916 -95 -37844
rect -45 -39916 -35 -37844
rect 1050 -37895 1120 -37705
rect 2160 -37756 2170 -35684
rect 2220 -37756 2230 -35684
rect 2160 -37844 2230 -37756
rect -105 -40004 -35 -39916
rect -1215 -42120 -1145 -42025
rect -105 -42076 -95 -40004
rect -45 -42076 -35 -40004
rect 1050 -40055 1120 -39865
rect 2160 -39916 2170 -37844
rect 2220 -39916 2230 -37844
rect 2160 -40004 2230 -39916
rect -105 -42120 -35 -42076
rect 1050 -42120 1120 -42025
rect 2160 -42076 2170 -40004
rect 2220 -42076 2230 -40004
rect 2160 -42120 2230 -42076
<< properties >>
string parameters w 20.00 l 20.00 val 413.6 carea 1.00 cperi 0.17 nx 2 ny 39 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
