magic
tech EFXH018D
timestamp 1523028597
<< metal1 >>
tri 3150 -225 3300 -75 se
rect 3300 -225 3450 75
tri 3000 -525 3150 -375 se
rect 3150 -525 3450 -225
rect 1650 -675 2250 -525
tri 1800 -825 1950 -675 ne
rect 1950 -825 2550 -675
rect 3000 -825 3300 -525
tri 3300 -675 3450 -525 nw
tri 3600 -675 3750 -525 se
rect 3750 -675 3900 -375
rect 1200 -1125 1800 -975
tri 1800 -1125 1950 -975 sw
tri 2100 -1125 2400 -825 ne
rect 2400 -975 3300 -825
rect 2400 -1125 2850 -975
tri 1350 -1275 1500 -1125 ne
rect 1500 -1275 2100 -1125
tri 2100 -1275 2250 -1125 sw
rect 750 -1575 1350 -1425
tri 1350 -1575 1500 -1425 sw
tri 1650 -1575 1950 -1275 ne
rect 1950 -1425 2400 -1275
tri 2400 -1425 2700 -1125 ne
rect 2700 -1425 2850 -1125
tri 2850 -1425 3300 -975 nw
tri 3450 -975 3600 -825 se
rect 3600 -975 3900 -675
tri 3300 -1275 3450 -1125 se
rect 3450 -1275 3750 -975
tri 3750 -1125 3900 -975 nw
tri 4050 -1125 4200 -975 se
rect 4200 -1125 4350 -825
rect 3300 -1425 3600 -1275
tri 3600 -1425 3750 -1275 nw
rect 1950 -1575 2250 -1425
tri 2250 -1575 2400 -1425 nw
tri 3300 -1575 3450 -1425 ne
rect 3450 -1575 3600 -1425
tri 3750 -1575 4050 -1275 se
rect 4050 -1425 4350 -1125
rect 4050 -1575 4200 -1425
tri 4200 -1575 4350 -1425 nw
tri 4500 -1575 4650 -1425 se
rect 4650 -1575 4800 -1275
tri 900 -1725 1050 -1575 ne
rect 1050 -1725 1650 -1575
tri 1650 -1725 1800 -1575 sw
rect 300 -2025 900 -1875
tri 900 -2025 1050 -1875 sw
tri 1200 -2025 1500 -1725 ne
rect 1500 -1875 1800 -1725
rect 3750 -1725 4200 -1575
tri 3750 -1875 3900 -1725 ne
rect 3900 -1875 4050 -1725
tri 4050 -1875 4200 -1725 nw
rect 1500 -2025 1650 -1875
tri 1650 -2025 1800 -1875 nw
tri 4200 -2025 4500 -1725 se
rect 4500 -1875 4800 -1575
rect 4500 -2025 4650 -1875
tri 4650 -2025 4800 -1875 nw
tri 5100 -1875 5250 -1725 se
rect 5250 -1875 5400 -1575
rect 5100 -2025 5400 -1875
tri 450 -2175 600 -2025 ne
rect 600 -2175 1350 -2025
tri 1350 -2175 1500 -2025 sw
rect 0 -2475 450 -2325
tri 450 -2475 600 -2325 sw
tri 750 -2475 1050 -2175 ne
rect 1050 -2325 1500 -2175
rect 1050 -2475 1350 -2325
tri 1350 -2475 1500 -2325 nw
rect 4200 -2175 4650 -2025
rect 4200 -2325 4500 -2175
tri 4500 -2325 4650 -2175 nw
tri 4200 -2475 4350 -2325 ne
rect 4350 -2475 4500 -2325
tri 4650 -2475 5100 -2025 se
rect 5100 -2475 5250 -2025
tri 5250 -2175 5400 -2025 nw
tri 150 -2775 450 -2475 ne
rect 450 -2775 900 -2475
tri 600 -2925 750 -2775 ne
rect 750 -2925 900 -2775
tri 900 -2925 1350 -2475 sw
tri 600 -3075 750 -2925 se
rect 750 -3075 1350 -2925
tri 450 -3375 600 -3225 se
rect 600 -3375 1050 -3075
tri 1050 -3375 1350 -3075 nw
tri 4350 -2775 4650 -2475 se
rect 4650 -2775 5100 -2475
tri 5100 -2625 5250 -2475 nw
rect 4350 -3075 4950 -2775
tri 4950 -2925 5100 -2775 nw
tri 4950 -3075 5100 -2925 sw
tri 4350 -3225 4500 -3075 ne
rect 4500 -3225 5250 -3075
tri 4650 -3375 4800 -3225 ne
rect 4800 -3375 5250 -3225
tri 5250 -3375 5550 -3075 sw
rect 450 -3675 750 -3375
tri 750 -3675 1050 -3375 nw
tri 1050 -3525 1200 -3375 se
rect 1200 -3525 1350 -3375
tri 1350 -3525 1500 -3375 sw
tri 300 -3825 450 -3675 se
rect 450 -3825 600 -3675
tri 600 -3825 750 -3675 nw
tri 900 -3825 1050 -3675 se
rect 1050 -3825 1500 -3525
tri 4200 -3525 4350 -3375 se
rect 4350 -3525 4500 -3375
rect 4200 -3675 4500 -3525
tri 4200 -3825 4350 -3675 ne
rect 4350 -3825 4500 -3675
tri 4500 -3825 4950 -3375 sw
tri 5100 -3525 5250 -3375 ne
rect 5250 -3525 5700 -3375
rect 300 -3975 600 -3825
rect 300 -4275 450 -3975
tri 450 -4125 600 -3975 nw
rect 900 -4125 1200 -3825
tri 1200 -4125 1500 -3825 nw
tri 1500 -3975 1650 -3825 se
rect 1650 -3975 1800 -3825
tri 1800 -3975 1950 -3825 sw
rect 1500 -4125 1950 -3975
tri 750 -4425 900 -4275 se
rect 900 -4425 1050 -4125
tri 1050 -4275 1200 -4125 nw
tri 1350 -4275 1500 -4125 se
rect 1500 -4275 1800 -4125
tri 1800 -4275 1950 -4125 nw
tri 3750 -3975 3900 -3825 se
rect 3900 -3975 4050 -3825
tri 4050 -3975 4200 -3825 sw
tri 4500 -3975 4650 -3825 ne
rect 4650 -3975 5250 -3825
rect 3750 -4125 4350 -3975
tri 3750 -4275 3900 -4125 ne
rect 3900 -4275 4350 -4125
tri 4350 -4275 4650 -3975 sw
rect 750 -4725 900 -4425
tri 900 -4575 1050 -4425 nw
rect 1350 -4425 1800 -4275
rect 1350 -5025 1500 -4425
tri 1500 -4725 1800 -4425 nw
tri 1950 -4425 2100 -4275 se
rect 2100 -4425 2250 -4275
tri 2250 -4425 2400 -4275 sw
tri 3300 -4425 3450 -4275 se
rect 3450 -4425 3600 -4275
tri 3600 -4425 3750 -4275 sw
tri 4050 -4425 4200 -4275 ne
rect 4200 -4425 4800 -4275
rect 1950 -4575 2400 -4425
tri 1800 -4725 1950 -4575 se
rect 1950 -4725 2100 -4575
rect 1800 -5025 2100 -4725
tri 2100 -4875 2400 -4575 nw
tri 2550 -4575 2700 -4425 se
rect 2700 -4575 3000 -4425
rect 2550 -4725 3000 -4575
tri 3000 -4725 3300 -4425 sw
rect 3300 -4575 3900 -4425
tri 3300 -4725 3450 -4575 ne
rect 3450 -4725 3900 -4575
tri 3900 -4725 4200 -4425 sw
tri 2400 -4875 2550 -4725 se
rect 2550 -4875 3300 -4725
rect 2400 -5025 3300 -4875
tri 3300 -5025 3600 -4725 sw
tri 3600 -4875 3750 -4725 ne
rect 3750 -4875 4500 -4725
rect 1800 -5325 1950 -5025
tri 1950 -5175 2100 -5025 nw
tri 2250 -5175 2400 -5025 se
rect 2400 -5175 2550 -5025
rect 2250 -5475 2550 -5175
tri 2550 -5325 2850 -5025 nw
tri 2850 -5175 3000 -5025 ne
rect 3000 -5175 3600 -5025
tri 3600 -5175 3750 -5025 sw
tri 3150 -5325 3300 -5175 ne
rect 3300 -5325 4050 -5175
rect 2250 -5775 2400 -5475
tri 2400 -5625 2550 -5475 nw
<< metal2 >>
tri 2550 -1875 2850 -1575 se
rect 2850 -1725 3300 -1575
tri 3300 -1725 3450 -1575 sw
rect 2850 -1875 3600 -1725
tri 3600 -1875 3750 -1725 sw
rect 2550 -2025 3750 -1875
rect 1950 -2175 2100 -2025
tri 2100 -2175 2250 -2025 sw
rect 2400 -2175 3750 -2025
tri 1650 -2625 1800 -2475 se
rect 1800 -2625 2250 -2175
rect 2550 -2325 3150 -2175
rect 3300 -2325 3600 -2175
rect 2550 -2475 3000 -2325
tri 3150 -2475 3300 -2325 se
rect 3300 -2475 3900 -2325
rect 2700 -2625 3900 -2475
tri 3900 -2625 4050 -2475 sw
rect 1650 -2775 1950 -2625
rect 2100 -2775 2250 -2625
rect 2850 -2775 4050 -2625
rect 1500 -2925 1950 -2775
rect 3150 -2925 4050 -2775
tri 4050 -2925 4200 -2775 sw
rect 1500 -3075 2250 -2925
rect 3150 -3075 3450 -2925
tri 3450 -3075 3600 -2925 nw
tri 3750 -3075 3900 -2925 ne
rect 3900 -3075 4200 -2925
rect 1500 -3225 1800 -3075
rect 1950 -3225 2250 -3075
tri 1500 -3375 1650 -3225 ne
rect 1650 -3525 2250 -3225
tri 2700 -3525 3000 -3225 se
rect 3000 -3375 3150 -3225
rect 3000 -3525 3300 -3375
rect 1650 -3675 2400 -3525
rect 2700 -3675 3300 -3525
tri 3300 -3675 3450 -3525 sw
tri 1650 -3825 1800 -3675 ne
rect 1800 -3825 2250 -3675
tri 2400 -3825 2550 -3675 se
rect 2550 -3825 3450 -3675
tri 1950 -3975 2100 -3825 ne
rect 2100 -3975 2400 -3825
tri 2400 -3975 2550 -3825 nw
rect 2700 -3975 3450 -3825
tri 3450 -3975 3600 -3825 sw
tri 3150 -4125 3300 -3975 ne
rect 3300 -4125 3600 -3975
<< end >>
