magic
tech EFXH018D
timestamp 1494891594
<< metal2 >>
rect 0 848 528 960
rect 0 528 104 848
rect 0 424 368 528
rect 0 104 104 424
rect 0 0 528 104
<< end >>
