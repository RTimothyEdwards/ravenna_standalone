magic
tech EFXH018D
magscale 1 2
timestamp 1565723183
<< mimcap >>
rect -79105 4130 -75105 4160
rect -79105 190 -79075 4130
rect -75135 190 -75105 4130
rect -79105 160 -75105 190
rect -74575 4130 -70575 4160
rect -74575 190 -74545 4130
rect -70605 190 -70575 4130
rect -74575 160 -70575 190
rect -70045 4130 -66045 4160
rect -70045 190 -70015 4130
rect -66075 190 -66045 4130
rect -70045 160 -66045 190
rect -65515 4130 -61515 4160
rect -65515 190 -65485 4130
rect -61545 190 -61515 4130
rect -65515 160 -61515 190
rect -60985 4130 -56985 4160
rect -60985 190 -60955 4130
rect -57015 190 -56985 4130
rect -60985 160 -56985 190
rect -56455 4130 -52455 4160
rect -56455 190 -56425 4130
rect -52485 190 -52455 4130
rect -56455 160 -52455 190
rect -51925 4130 -47925 4160
rect -51925 190 -51895 4130
rect -47955 190 -47925 4130
rect -51925 160 -47925 190
rect -47395 4130 -43395 4160
rect -47395 190 -47365 4130
rect -43425 190 -43395 4130
rect -47395 160 -43395 190
rect -42865 4130 -38865 4160
rect -42865 190 -42835 4130
rect -38895 190 -38865 4130
rect -42865 160 -38865 190
rect -38335 4130 -34335 4160
rect -38335 190 -38305 4130
rect -34365 190 -34335 4130
rect -38335 160 -34335 190
rect -33805 4130 -29805 4160
rect -33805 190 -33775 4130
rect -29835 190 -29805 4130
rect -33805 160 -29805 190
rect -29275 4130 -25275 4160
rect -29275 190 -29245 4130
rect -25305 190 -25275 4130
rect -29275 160 -25275 190
rect -24745 4130 -20745 4160
rect -24745 190 -24715 4130
rect -20775 190 -20745 4130
rect -24745 160 -20745 190
rect -20215 4130 -16215 4160
rect -20215 190 -20185 4130
rect -16245 190 -16215 4130
rect -20215 160 -16215 190
rect -15685 4130 -11685 4160
rect -15685 190 -15655 4130
rect -11715 190 -11685 4130
rect -15685 160 -11685 190
rect -11155 4130 -7155 4160
rect -11155 190 -11125 4130
rect -7185 190 -7155 4130
rect -11155 160 -7155 190
rect -6625 4130 -2625 4160
rect -6625 190 -6595 4130
rect -2655 190 -2625 4130
rect -6625 160 -2625 190
rect -2095 4130 1905 4160
rect -2095 190 -2065 4130
rect 1875 190 1905 4130
rect -2095 160 1905 190
rect 2435 4130 6435 4160
rect 2435 190 2465 4130
rect 6405 190 6435 4130
rect 2435 160 6435 190
rect 6965 4130 10965 4160
rect 6965 190 6995 4130
rect 10935 190 10965 4130
rect 6965 160 10965 190
rect 11495 4130 15495 4160
rect 11495 190 11525 4130
rect 15465 190 15495 4130
rect 11495 160 15495 190
rect 16025 4130 20025 4160
rect 16025 190 16055 4130
rect 19995 190 20025 4130
rect 16025 160 20025 190
rect 20555 4130 24555 4160
rect 20555 190 20585 4130
rect 24525 190 24555 4130
rect 20555 160 24555 190
rect 25085 4130 29085 4160
rect 25085 190 25115 4130
rect 29055 190 29085 4130
rect 25085 160 29085 190
rect 29615 4130 33615 4160
rect 29615 190 29645 4130
rect 33585 190 33615 4130
rect 29615 160 33615 190
rect 34145 4130 38145 4160
rect 34145 190 34175 4130
rect 38115 190 38145 4130
rect 34145 160 38145 190
rect 38675 4130 42675 4160
rect 38675 190 38705 4130
rect 42645 190 42675 4130
rect 38675 160 42675 190
rect 43205 4130 47205 4160
rect 43205 190 43235 4130
rect 47175 190 47205 4130
rect 43205 160 47205 190
rect 47735 4130 51735 4160
rect 47735 190 47765 4130
rect 51705 190 51735 4130
rect 47735 160 51735 190
rect 52265 4130 56265 4160
rect 52265 190 52295 4130
rect 56235 190 56265 4130
rect 52265 160 56265 190
rect 56795 4130 60795 4160
rect 56795 190 56825 4130
rect 60765 190 60795 4130
rect 56795 160 60795 190
rect 61325 4130 65325 4160
rect 61325 190 61355 4130
rect 65295 190 65325 4130
rect 61325 160 65325 190
rect 65855 4130 69855 4160
rect 65855 190 65885 4130
rect 69825 190 69855 4130
rect 65855 160 69855 190
rect 70385 4130 74385 4160
rect 70385 190 70415 4130
rect 74355 190 74385 4130
rect 70385 160 74385 190
rect 74915 4130 78915 4160
rect 74915 190 74945 4130
rect 78885 190 78915 4130
rect 74915 160 78915 190
rect -79105 -190 -75105 -160
rect -79105 -4130 -79075 -190
rect -75135 -4130 -75105 -190
rect -79105 -4160 -75105 -4130
rect -74575 -190 -70575 -160
rect -74575 -4130 -74545 -190
rect -70605 -4130 -70575 -190
rect -74575 -4160 -70575 -4130
rect -70045 -190 -66045 -160
rect -70045 -4130 -70015 -190
rect -66075 -4130 -66045 -190
rect -70045 -4160 -66045 -4130
rect -65515 -190 -61515 -160
rect -65515 -4130 -65485 -190
rect -61545 -4130 -61515 -190
rect -65515 -4160 -61515 -4130
rect -60985 -190 -56985 -160
rect -60985 -4130 -60955 -190
rect -57015 -4130 -56985 -190
rect -60985 -4160 -56985 -4130
rect -56455 -190 -52455 -160
rect -56455 -4130 -56425 -190
rect -52485 -4130 -52455 -190
rect -56455 -4160 -52455 -4130
rect -51925 -190 -47925 -160
rect -51925 -4130 -51895 -190
rect -47955 -4130 -47925 -190
rect -51925 -4160 -47925 -4130
rect -47395 -190 -43395 -160
rect -47395 -4130 -47365 -190
rect -43425 -4130 -43395 -190
rect -47395 -4160 -43395 -4130
rect -42865 -190 -38865 -160
rect -42865 -4130 -42835 -190
rect -38895 -4130 -38865 -190
rect -42865 -4160 -38865 -4130
rect -38335 -190 -34335 -160
rect -38335 -4130 -38305 -190
rect -34365 -4130 -34335 -190
rect -38335 -4160 -34335 -4130
rect -33805 -190 -29805 -160
rect -33805 -4130 -33775 -190
rect -29835 -4130 -29805 -190
rect -33805 -4160 -29805 -4130
rect -29275 -190 -25275 -160
rect -29275 -4130 -29245 -190
rect -25305 -4130 -25275 -190
rect -29275 -4160 -25275 -4130
rect -24745 -190 -20745 -160
rect -24745 -4130 -24715 -190
rect -20775 -4130 -20745 -190
rect -24745 -4160 -20745 -4130
rect -20215 -190 -16215 -160
rect -20215 -4130 -20185 -190
rect -16245 -4130 -16215 -190
rect -20215 -4160 -16215 -4130
rect -15685 -190 -11685 -160
rect -15685 -4130 -15655 -190
rect -11715 -4130 -11685 -190
rect -15685 -4160 -11685 -4130
rect -11155 -190 -7155 -160
rect -11155 -4130 -11125 -190
rect -7185 -4130 -7155 -190
rect -11155 -4160 -7155 -4130
rect -6625 -190 -2625 -160
rect -6625 -4130 -6595 -190
rect -2655 -4130 -2625 -190
rect -6625 -4160 -2625 -4130
rect -2095 -190 1905 -160
rect -2095 -4130 -2065 -190
rect 1875 -4130 1905 -190
rect -2095 -4160 1905 -4130
rect 2435 -190 6435 -160
rect 2435 -4130 2465 -190
rect 6405 -4130 6435 -190
rect 2435 -4160 6435 -4130
rect 6965 -190 10965 -160
rect 6965 -4130 6995 -190
rect 10935 -4130 10965 -190
rect 6965 -4160 10965 -4130
rect 11495 -190 15495 -160
rect 11495 -4130 11525 -190
rect 15465 -4130 15495 -190
rect 11495 -4160 15495 -4130
rect 16025 -190 20025 -160
rect 16025 -4130 16055 -190
rect 19995 -4130 20025 -190
rect 16025 -4160 20025 -4130
rect 20555 -190 24555 -160
rect 20555 -4130 20585 -190
rect 24525 -4130 24555 -190
rect 20555 -4160 24555 -4130
rect 25085 -190 29085 -160
rect 25085 -4130 25115 -190
rect 29055 -4130 29085 -190
rect 25085 -4160 29085 -4130
rect 29615 -190 33615 -160
rect 29615 -4130 29645 -190
rect 33585 -4130 33615 -190
rect 29615 -4160 33615 -4130
rect 34145 -190 38145 -160
rect 34145 -4130 34175 -190
rect 38115 -4130 38145 -190
rect 34145 -4160 38145 -4130
rect 38675 -190 42675 -160
rect 38675 -4130 38705 -190
rect 42645 -4130 42675 -190
rect 38675 -4160 42675 -4130
rect 43205 -190 47205 -160
rect 43205 -4130 43235 -190
rect 47175 -4130 47205 -190
rect 43205 -4160 47205 -4130
rect 47735 -190 51735 -160
rect 47735 -4130 47765 -190
rect 51705 -4130 51735 -190
rect 47735 -4160 51735 -4130
rect 52265 -190 56265 -160
rect 52265 -4130 52295 -190
rect 56235 -4130 56265 -190
rect 52265 -4160 56265 -4130
rect 56795 -190 60795 -160
rect 56795 -4130 56825 -190
rect 60765 -4130 60795 -190
rect 56795 -4160 60795 -4130
rect 61325 -190 65325 -160
rect 61325 -4130 61355 -190
rect 65295 -4130 65325 -190
rect 61325 -4160 65325 -4130
rect 65855 -190 69855 -160
rect 65855 -4130 65885 -190
rect 69825 -4130 69855 -190
rect 65855 -4160 69855 -4130
rect 70385 -190 74385 -160
rect 70385 -4130 70415 -190
rect 74355 -4130 74385 -190
rect 70385 -4160 74385 -4130
rect 74915 -190 78915 -160
rect 74915 -4130 74945 -190
rect 78885 -4130 78915 -190
rect 74915 -4160 78915 -4130
<< mimcapcontact >>
rect -79075 190 -75135 4130
rect -74545 190 -70605 4130
rect -70015 190 -66075 4130
rect -65485 190 -61545 4130
rect -60955 190 -57015 4130
rect -56425 190 -52485 4130
rect -51895 190 -47955 4130
rect -47365 190 -43425 4130
rect -42835 190 -38895 4130
rect -38305 190 -34365 4130
rect -33775 190 -29835 4130
rect -29245 190 -25305 4130
rect -24715 190 -20775 4130
rect -20185 190 -16245 4130
rect -15655 190 -11715 4130
rect -11125 190 -7185 4130
rect -6595 190 -2655 4130
rect -2065 190 1875 4130
rect 2465 190 6405 4130
rect 6995 190 10935 4130
rect 11525 190 15465 4130
rect 16055 190 19995 4130
rect 20585 190 24525 4130
rect 25115 190 29055 4130
rect 29645 190 33585 4130
rect 34175 190 38115 4130
rect 38705 190 42645 4130
rect 43235 190 47175 4130
rect 47765 190 51705 4130
rect 52295 190 56235 4130
rect 56825 190 60765 4130
rect 61355 190 65295 4130
rect 65885 190 69825 4130
rect 70415 190 74355 4130
rect 74945 190 78885 4130
rect -79075 -4130 -75135 -190
rect -74545 -4130 -70605 -190
rect -70015 -4130 -66075 -190
rect -65485 -4130 -61545 -190
rect -60955 -4130 -57015 -190
rect -56425 -4130 -52485 -190
rect -51895 -4130 -47955 -190
rect -47365 -4130 -43425 -190
rect -42835 -4130 -38895 -190
rect -38305 -4130 -34365 -190
rect -33775 -4130 -29835 -190
rect -29245 -4130 -25305 -190
rect -24715 -4130 -20775 -190
rect -20185 -4130 -16245 -190
rect -15655 -4130 -11715 -190
rect -11125 -4130 -7185 -190
rect -6595 -4130 -2655 -190
rect -2065 -4130 1875 -190
rect 2465 -4130 6405 -190
rect 6995 -4130 10935 -190
rect 11525 -4130 15465 -190
rect 16055 -4130 19995 -190
rect 20585 -4130 24525 -190
rect 25115 -4130 29055 -190
rect 29645 -4130 33585 -190
rect 34175 -4130 38115 -190
rect 38705 -4130 42645 -190
rect 43235 -4130 47175 -190
rect 47765 -4130 51705 -190
rect 52295 -4130 56235 -190
rect 56825 -4130 60765 -190
rect 61355 -4130 65295 -190
rect 65885 -4130 69825 -190
rect 70415 -4130 74355 -190
rect 74945 -4130 78885 -190
<< metal4 >>
rect -79205 4232 -74815 4260
rect -79205 4160 -74935 4232
rect -79205 160 -79105 4160
rect -75105 160 -74935 4160
rect -79205 88 -74935 160
rect -74835 88 -74815 4232
rect -79205 60 -74815 88
rect -74675 4232 -70285 4260
rect -74675 4160 -70405 4232
rect -74675 160 -74575 4160
rect -70575 160 -70405 4160
rect -74675 88 -70405 160
rect -70305 88 -70285 4232
rect -74675 60 -70285 88
rect -70145 4232 -65755 4260
rect -70145 4160 -65875 4232
rect -70145 160 -70045 4160
rect -66045 160 -65875 4160
rect -70145 88 -65875 160
rect -65775 88 -65755 4232
rect -70145 60 -65755 88
rect -65615 4232 -61225 4260
rect -65615 4160 -61345 4232
rect -65615 160 -65515 4160
rect -61515 160 -61345 4160
rect -65615 88 -61345 160
rect -61245 88 -61225 4232
rect -65615 60 -61225 88
rect -61085 4232 -56695 4260
rect -61085 4160 -56815 4232
rect -61085 160 -60985 4160
rect -56985 160 -56815 4160
rect -61085 88 -56815 160
rect -56715 88 -56695 4232
rect -61085 60 -56695 88
rect -56555 4232 -52165 4260
rect -56555 4160 -52285 4232
rect -56555 160 -56455 4160
rect -52455 160 -52285 4160
rect -56555 88 -52285 160
rect -52185 88 -52165 4232
rect -56555 60 -52165 88
rect -52025 4232 -47635 4260
rect -52025 4160 -47755 4232
rect -52025 160 -51925 4160
rect -47925 160 -47755 4160
rect -52025 88 -47755 160
rect -47655 88 -47635 4232
rect -52025 60 -47635 88
rect -47495 4232 -43105 4260
rect -47495 4160 -43225 4232
rect -47495 160 -47395 4160
rect -43395 160 -43225 4160
rect -47495 88 -43225 160
rect -43125 88 -43105 4232
rect -47495 60 -43105 88
rect -42965 4232 -38575 4260
rect -42965 4160 -38695 4232
rect -42965 160 -42865 4160
rect -38865 160 -38695 4160
rect -42965 88 -38695 160
rect -38595 88 -38575 4232
rect -42965 60 -38575 88
rect -38435 4232 -34045 4260
rect -38435 4160 -34165 4232
rect -38435 160 -38335 4160
rect -34335 160 -34165 4160
rect -38435 88 -34165 160
rect -34065 88 -34045 4232
rect -38435 60 -34045 88
rect -33905 4232 -29515 4260
rect -33905 4160 -29635 4232
rect -33905 160 -33805 4160
rect -29805 160 -29635 4160
rect -33905 88 -29635 160
rect -29535 88 -29515 4232
rect -33905 60 -29515 88
rect -29375 4232 -24985 4260
rect -29375 4160 -25105 4232
rect -29375 160 -29275 4160
rect -25275 160 -25105 4160
rect -29375 88 -25105 160
rect -25005 88 -24985 4232
rect -29375 60 -24985 88
rect -24845 4232 -20455 4260
rect -24845 4160 -20575 4232
rect -24845 160 -24745 4160
rect -20745 160 -20575 4160
rect -24845 88 -20575 160
rect -20475 88 -20455 4232
rect -24845 60 -20455 88
rect -20315 4232 -15925 4260
rect -20315 4160 -16045 4232
rect -20315 160 -20215 4160
rect -16215 160 -16045 4160
rect -20315 88 -16045 160
rect -15945 88 -15925 4232
rect -20315 60 -15925 88
rect -15785 4232 -11395 4260
rect -15785 4160 -11515 4232
rect -15785 160 -15685 4160
rect -11685 160 -11515 4160
rect -15785 88 -11515 160
rect -11415 88 -11395 4232
rect -15785 60 -11395 88
rect -11255 4232 -6865 4260
rect -11255 4160 -6985 4232
rect -11255 160 -11155 4160
rect -7155 160 -6985 4160
rect -11255 88 -6985 160
rect -6885 88 -6865 4232
rect -11255 60 -6865 88
rect -6725 4232 -2335 4260
rect -6725 4160 -2455 4232
rect -6725 160 -6625 4160
rect -2625 160 -2455 4160
rect -6725 88 -2455 160
rect -2355 88 -2335 4232
rect -6725 60 -2335 88
rect -2195 4232 2195 4260
rect -2195 4160 2075 4232
rect -2195 160 -2095 4160
rect 1905 160 2075 4160
rect -2195 88 2075 160
rect 2175 88 2195 4232
rect -2195 60 2195 88
rect 2335 4232 6725 4260
rect 2335 4160 6605 4232
rect 2335 160 2435 4160
rect 6435 160 6605 4160
rect 2335 88 6605 160
rect 6705 88 6725 4232
rect 2335 60 6725 88
rect 6865 4232 11255 4260
rect 6865 4160 11135 4232
rect 6865 160 6965 4160
rect 10965 160 11135 4160
rect 6865 88 11135 160
rect 11235 88 11255 4232
rect 6865 60 11255 88
rect 11395 4232 15785 4260
rect 11395 4160 15665 4232
rect 11395 160 11495 4160
rect 15495 160 15665 4160
rect 11395 88 15665 160
rect 15765 88 15785 4232
rect 11395 60 15785 88
rect 15925 4232 20315 4260
rect 15925 4160 20195 4232
rect 15925 160 16025 4160
rect 20025 160 20195 4160
rect 15925 88 20195 160
rect 20295 88 20315 4232
rect 15925 60 20315 88
rect 20455 4232 24845 4260
rect 20455 4160 24725 4232
rect 20455 160 20555 4160
rect 24555 160 24725 4160
rect 20455 88 24725 160
rect 24825 88 24845 4232
rect 20455 60 24845 88
rect 24985 4232 29375 4260
rect 24985 4160 29255 4232
rect 24985 160 25085 4160
rect 29085 160 29255 4160
rect 24985 88 29255 160
rect 29355 88 29375 4232
rect 24985 60 29375 88
rect 29515 4232 33905 4260
rect 29515 4160 33785 4232
rect 29515 160 29615 4160
rect 33615 160 33785 4160
rect 29515 88 33785 160
rect 33885 88 33905 4232
rect 29515 60 33905 88
rect 34045 4232 38435 4260
rect 34045 4160 38315 4232
rect 34045 160 34145 4160
rect 38145 160 38315 4160
rect 34045 88 38315 160
rect 38415 88 38435 4232
rect 34045 60 38435 88
rect 38575 4232 42965 4260
rect 38575 4160 42845 4232
rect 38575 160 38675 4160
rect 42675 160 42845 4160
rect 38575 88 42845 160
rect 42945 88 42965 4232
rect 38575 60 42965 88
rect 43105 4232 47495 4260
rect 43105 4160 47375 4232
rect 43105 160 43205 4160
rect 47205 160 47375 4160
rect 43105 88 47375 160
rect 47475 88 47495 4232
rect 43105 60 47495 88
rect 47635 4232 52025 4260
rect 47635 4160 51905 4232
rect 47635 160 47735 4160
rect 51735 160 51905 4160
rect 47635 88 51905 160
rect 52005 88 52025 4232
rect 47635 60 52025 88
rect 52165 4232 56555 4260
rect 52165 4160 56435 4232
rect 52165 160 52265 4160
rect 56265 160 56435 4160
rect 52165 88 56435 160
rect 56535 88 56555 4232
rect 52165 60 56555 88
rect 56695 4232 61085 4260
rect 56695 4160 60965 4232
rect 56695 160 56795 4160
rect 60795 160 60965 4160
rect 56695 88 60965 160
rect 61065 88 61085 4232
rect 56695 60 61085 88
rect 61225 4232 65615 4260
rect 61225 4160 65495 4232
rect 61225 160 61325 4160
rect 65325 160 65495 4160
rect 61225 88 65495 160
rect 65595 88 65615 4232
rect 61225 60 65615 88
rect 65755 4232 70145 4260
rect 65755 4160 70025 4232
rect 65755 160 65855 4160
rect 69855 160 70025 4160
rect 65755 88 70025 160
rect 70125 88 70145 4232
rect 65755 60 70145 88
rect 70285 4232 74675 4260
rect 70285 4160 74555 4232
rect 70285 160 70385 4160
rect 74385 160 74555 4160
rect 70285 88 74555 160
rect 74655 88 74675 4232
rect 70285 60 74675 88
rect 74815 4232 79205 4260
rect 74815 4160 79085 4232
rect 74815 160 74915 4160
rect 78915 160 79085 4160
rect 74815 88 79085 160
rect 79185 88 79205 4232
rect 74815 60 79205 88
rect -79205 -88 -74815 -60
rect -79205 -160 -74935 -88
rect -79205 -4160 -79105 -160
rect -75105 -4160 -74935 -160
rect -79205 -4232 -74935 -4160
rect -74835 -4232 -74815 -88
rect -79205 -4260 -74815 -4232
rect -74675 -88 -70285 -60
rect -74675 -160 -70405 -88
rect -74675 -4160 -74575 -160
rect -70575 -4160 -70405 -160
rect -74675 -4232 -70405 -4160
rect -70305 -4232 -70285 -88
rect -74675 -4260 -70285 -4232
rect -70145 -88 -65755 -60
rect -70145 -160 -65875 -88
rect -70145 -4160 -70045 -160
rect -66045 -4160 -65875 -160
rect -70145 -4232 -65875 -4160
rect -65775 -4232 -65755 -88
rect -70145 -4260 -65755 -4232
rect -65615 -88 -61225 -60
rect -65615 -160 -61345 -88
rect -65615 -4160 -65515 -160
rect -61515 -4160 -61345 -160
rect -65615 -4232 -61345 -4160
rect -61245 -4232 -61225 -88
rect -65615 -4260 -61225 -4232
rect -61085 -88 -56695 -60
rect -61085 -160 -56815 -88
rect -61085 -4160 -60985 -160
rect -56985 -4160 -56815 -160
rect -61085 -4232 -56815 -4160
rect -56715 -4232 -56695 -88
rect -61085 -4260 -56695 -4232
rect -56555 -88 -52165 -60
rect -56555 -160 -52285 -88
rect -56555 -4160 -56455 -160
rect -52455 -4160 -52285 -160
rect -56555 -4232 -52285 -4160
rect -52185 -4232 -52165 -88
rect -56555 -4260 -52165 -4232
rect -52025 -88 -47635 -60
rect -52025 -160 -47755 -88
rect -52025 -4160 -51925 -160
rect -47925 -4160 -47755 -160
rect -52025 -4232 -47755 -4160
rect -47655 -4232 -47635 -88
rect -52025 -4260 -47635 -4232
rect -47495 -88 -43105 -60
rect -47495 -160 -43225 -88
rect -47495 -4160 -47395 -160
rect -43395 -4160 -43225 -160
rect -47495 -4232 -43225 -4160
rect -43125 -4232 -43105 -88
rect -47495 -4260 -43105 -4232
rect -42965 -88 -38575 -60
rect -42965 -160 -38695 -88
rect -42965 -4160 -42865 -160
rect -38865 -4160 -38695 -160
rect -42965 -4232 -38695 -4160
rect -38595 -4232 -38575 -88
rect -42965 -4260 -38575 -4232
rect -38435 -88 -34045 -60
rect -38435 -160 -34165 -88
rect -38435 -4160 -38335 -160
rect -34335 -4160 -34165 -160
rect -38435 -4232 -34165 -4160
rect -34065 -4232 -34045 -88
rect -38435 -4260 -34045 -4232
rect -33905 -88 -29515 -60
rect -33905 -160 -29635 -88
rect -33905 -4160 -33805 -160
rect -29805 -4160 -29635 -160
rect -33905 -4232 -29635 -4160
rect -29535 -4232 -29515 -88
rect -33905 -4260 -29515 -4232
rect -29375 -88 -24985 -60
rect -29375 -160 -25105 -88
rect -29375 -4160 -29275 -160
rect -25275 -4160 -25105 -160
rect -29375 -4232 -25105 -4160
rect -25005 -4232 -24985 -88
rect -29375 -4260 -24985 -4232
rect -24845 -88 -20455 -60
rect -24845 -160 -20575 -88
rect -24845 -4160 -24745 -160
rect -20745 -4160 -20575 -160
rect -24845 -4232 -20575 -4160
rect -20475 -4232 -20455 -88
rect -24845 -4260 -20455 -4232
rect -20315 -88 -15925 -60
rect -20315 -160 -16045 -88
rect -20315 -4160 -20215 -160
rect -16215 -4160 -16045 -160
rect -20315 -4232 -16045 -4160
rect -15945 -4232 -15925 -88
rect -20315 -4260 -15925 -4232
rect -15785 -88 -11395 -60
rect -15785 -160 -11515 -88
rect -15785 -4160 -15685 -160
rect -11685 -4160 -11515 -160
rect -15785 -4232 -11515 -4160
rect -11415 -4232 -11395 -88
rect -15785 -4260 -11395 -4232
rect -11255 -88 -6865 -60
rect -11255 -160 -6985 -88
rect -11255 -4160 -11155 -160
rect -7155 -4160 -6985 -160
rect -11255 -4232 -6985 -4160
rect -6885 -4232 -6865 -88
rect -11255 -4260 -6865 -4232
rect -6725 -88 -2335 -60
rect -6725 -160 -2455 -88
rect -6725 -4160 -6625 -160
rect -2625 -4160 -2455 -160
rect -6725 -4232 -2455 -4160
rect -2355 -4232 -2335 -88
rect -6725 -4260 -2335 -4232
rect -2195 -88 2195 -60
rect -2195 -160 2075 -88
rect -2195 -4160 -2095 -160
rect 1905 -4160 2075 -160
rect -2195 -4232 2075 -4160
rect 2175 -4232 2195 -88
rect -2195 -4260 2195 -4232
rect 2335 -88 6725 -60
rect 2335 -160 6605 -88
rect 2335 -4160 2435 -160
rect 6435 -4160 6605 -160
rect 2335 -4232 6605 -4160
rect 6705 -4232 6725 -88
rect 2335 -4260 6725 -4232
rect 6865 -88 11255 -60
rect 6865 -160 11135 -88
rect 6865 -4160 6965 -160
rect 10965 -4160 11135 -160
rect 6865 -4232 11135 -4160
rect 11235 -4232 11255 -88
rect 6865 -4260 11255 -4232
rect 11395 -88 15785 -60
rect 11395 -160 15665 -88
rect 11395 -4160 11495 -160
rect 15495 -4160 15665 -160
rect 11395 -4232 15665 -4160
rect 15765 -4232 15785 -88
rect 11395 -4260 15785 -4232
rect 15925 -88 20315 -60
rect 15925 -160 20195 -88
rect 15925 -4160 16025 -160
rect 20025 -4160 20195 -160
rect 15925 -4232 20195 -4160
rect 20295 -4232 20315 -88
rect 15925 -4260 20315 -4232
rect 20455 -88 24845 -60
rect 20455 -160 24725 -88
rect 20455 -4160 20555 -160
rect 24555 -4160 24725 -160
rect 20455 -4232 24725 -4160
rect 24825 -4232 24845 -88
rect 20455 -4260 24845 -4232
rect 24985 -88 29375 -60
rect 24985 -160 29255 -88
rect 24985 -4160 25085 -160
rect 29085 -4160 29255 -160
rect 24985 -4232 29255 -4160
rect 29355 -4232 29375 -88
rect 24985 -4260 29375 -4232
rect 29515 -88 33905 -60
rect 29515 -160 33785 -88
rect 29515 -4160 29615 -160
rect 33615 -4160 33785 -160
rect 29515 -4232 33785 -4160
rect 33885 -4232 33905 -88
rect 29515 -4260 33905 -4232
rect 34045 -88 38435 -60
rect 34045 -160 38315 -88
rect 34045 -4160 34145 -160
rect 38145 -4160 38315 -160
rect 34045 -4232 38315 -4160
rect 38415 -4232 38435 -88
rect 34045 -4260 38435 -4232
rect 38575 -88 42965 -60
rect 38575 -160 42845 -88
rect 38575 -4160 38675 -160
rect 42675 -4160 42845 -160
rect 38575 -4232 42845 -4160
rect 42945 -4232 42965 -88
rect 38575 -4260 42965 -4232
rect 43105 -88 47495 -60
rect 43105 -160 47375 -88
rect 43105 -4160 43205 -160
rect 47205 -4160 47375 -160
rect 43105 -4232 47375 -4160
rect 47475 -4232 47495 -88
rect 43105 -4260 47495 -4232
rect 47635 -88 52025 -60
rect 47635 -160 51905 -88
rect 47635 -4160 47735 -160
rect 51735 -4160 51905 -160
rect 47635 -4232 51905 -4160
rect 52005 -4232 52025 -88
rect 47635 -4260 52025 -4232
rect 52165 -88 56555 -60
rect 52165 -160 56435 -88
rect 52165 -4160 52265 -160
rect 56265 -4160 56435 -160
rect 52165 -4232 56435 -4160
rect 56535 -4232 56555 -88
rect 52165 -4260 56555 -4232
rect 56695 -88 61085 -60
rect 56695 -160 60965 -88
rect 56695 -4160 56795 -160
rect 60795 -4160 60965 -160
rect 56695 -4232 60965 -4160
rect 61065 -4232 61085 -88
rect 56695 -4260 61085 -4232
rect 61225 -88 65615 -60
rect 61225 -160 65495 -88
rect 61225 -4160 61325 -160
rect 65325 -4160 65495 -160
rect 61225 -4232 65495 -4160
rect 65595 -4232 65615 -88
rect 61225 -4260 65615 -4232
rect 65755 -88 70145 -60
rect 65755 -160 70025 -88
rect 65755 -4160 65855 -160
rect 69855 -4160 70025 -160
rect 65755 -4232 70025 -4160
rect 70125 -4232 70145 -88
rect 65755 -4260 70145 -4232
rect 70285 -88 74675 -60
rect 70285 -160 74555 -88
rect 70285 -4160 70385 -160
rect 74385 -4160 74555 -160
rect 70285 -4232 74555 -4160
rect 74655 -4232 74675 -88
rect 70285 -4260 74675 -4232
rect 74815 -88 79205 -60
rect 74815 -160 79085 -88
rect 74815 -4160 74915 -160
rect 78915 -4160 79085 -160
rect 74815 -4232 79085 -4160
rect 79185 -4232 79205 -88
rect 74815 -4260 79205 -4232
<< viatp >>
rect -74935 88 -74835 4232
rect -70405 88 -70305 4232
rect -65875 88 -65775 4232
rect -61345 88 -61245 4232
rect -56815 88 -56715 4232
rect -52285 88 -52185 4232
rect -47755 88 -47655 4232
rect -43225 88 -43125 4232
rect -38695 88 -38595 4232
rect -34165 88 -34065 4232
rect -29635 88 -29535 4232
rect -25105 88 -25005 4232
rect -20575 88 -20475 4232
rect -16045 88 -15945 4232
rect -11515 88 -11415 4232
rect -6985 88 -6885 4232
rect -2455 88 -2355 4232
rect 2075 88 2175 4232
rect 6605 88 6705 4232
rect 11135 88 11235 4232
rect 15665 88 15765 4232
rect 20195 88 20295 4232
rect 24725 88 24825 4232
rect 29255 88 29355 4232
rect 33785 88 33885 4232
rect 38315 88 38415 4232
rect 42845 88 42945 4232
rect 47375 88 47475 4232
rect 51905 88 52005 4232
rect 56435 88 56535 4232
rect 60965 88 61065 4232
rect 65495 88 65595 4232
rect 70025 88 70125 4232
rect 74555 88 74655 4232
rect 79085 88 79185 4232
rect -74935 -4232 -74835 -88
rect -70405 -4232 -70305 -88
rect -65875 -4232 -65775 -88
rect -61345 -4232 -61245 -88
rect -56815 -4232 -56715 -88
rect -52285 -4232 -52185 -88
rect -47755 -4232 -47655 -88
rect -43225 -4232 -43125 -88
rect -38695 -4232 -38595 -88
rect -34165 -4232 -34065 -88
rect -29635 -4232 -29535 -88
rect -25105 -4232 -25005 -88
rect -20575 -4232 -20475 -88
rect -16045 -4232 -15945 -88
rect -11515 -4232 -11415 -88
rect -6985 -4232 -6885 -88
rect -2455 -4232 -2355 -88
rect 2075 -4232 2175 -88
rect 6605 -4232 6705 -88
rect 11135 -4232 11235 -88
rect 15665 -4232 15765 -88
rect 20195 -4232 20295 -88
rect 24725 -4232 24825 -88
rect 29255 -4232 29355 -88
rect 33785 -4232 33885 -88
rect 38315 -4232 38415 -88
rect 42845 -4232 42945 -88
rect 47375 -4232 47475 -88
rect 51905 -4232 52005 -88
rect 56435 -4232 56535 -88
rect 60965 -4232 61065 -88
rect 65495 -4232 65595 -88
rect 70025 -4232 70125 -88
rect 74555 -4232 74655 -88
rect 79085 -4232 79185 -88
<< metaltp >>
rect -77175 4130 -77035 4320
rect -74955 4232 -74815 4320
rect -77175 -190 -77035 190
rect -74955 88 -74935 4232
rect -74835 88 -74815 4232
rect -72645 4130 -72505 4320
rect -70425 4232 -70285 4320
rect -74955 -88 -74815 88
rect -77175 -4320 -77035 -4130
rect -74955 -4232 -74935 -88
rect -74835 -4232 -74815 -88
rect -72645 -190 -72505 190
rect -70425 88 -70405 4232
rect -70305 88 -70285 4232
rect -68115 4130 -67975 4320
rect -65895 4232 -65755 4320
rect -70425 -88 -70285 88
rect -74955 -4320 -74815 -4232
rect -72645 -4320 -72505 -4130
rect -70425 -4232 -70405 -88
rect -70305 -4232 -70285 -88
rect -68115 -190 -67975 190
rect -65895 88 -65875 4232
rect -65775 88 -65755 4232
rect -63585 4130 -63445 4320
rect -61365 4232 -61225 4320
rect -65895 -88 -65755 88
rect -70425 -4320 -70285 -4232
rect -68115 -4320 -67975 -4130
rect -65895 -4232 -65875 -88
rect -65775 -4232 -65755 -88
rect -63585 -190 -63445 190
rect -61365 88 -61345 4232
rect -61245 88 -61225 4232
rect -59055 4130 -58915 4320
rect -56835 4232 -56695 4320
rect -61365 -88 -61225 88
rect -65895 -4320 -65755 -4232
rect -63585 -4320 -63445 -4130
rect -61365 -4232 -61345 -88
rect -61245 -4232 -61225 -88
rect -59055 -190 -58915 190
rect -56835 88 -56815 4232
rect -56715 88 -56695 4232
rect -54525 4130 -54385 4320
rect -52305 4232 -52165 4320
rect -56835 -88 -56695 88
rect -61365 -4320 -61225 -4232
rect -59055 -4320 -58915 -4130
rect -56835 -4232 -56815 -88
rect -56715 -4232 -56695 -88
rect -54525 -190 -54385 190
rect -52305 88 -52285 4232
rect -52185 88 -52165 4232
rect -49995 4130 -49855 4320
rect -47775 4232 -47635 4320
rect -52305 -88 -52165 88
rect -56835 -4320 -56695 -4232
rect -54525 -4320 -54385 -4130
rect -52305 -4232 -52285 -88
rect -52185 -4232 -52165 -88
rect -49995 -190 -49855 190
rect -47775 88 -47755 4232
rect -47655 88 -47635 4232
rect -45465 4130 -45325 4320
rect -43245 4232 -43105 4320
rect -47775 -88 -47635 88
rect -52305 -4320 -52165 -4232
rect -49995 -4320 -49855 -4130
rect -47775 -4232 -47755 -88
rect -47655 -4232 -47635 -88
rect -45465 -190 -45325 190
rect -43245 88 -43225 4232
rect -43125 88 -43105 4232
rect -40935 4130 -40795 4320
rect -38715 4232 -38575 4320
rect -43245 -88 -43105 88
rect -47775 -4320 -47635 -4232
rect -45465 -4320 -45325 -4130
rect -43245 -4232 -43225 -88
rect -43125 -4232 -43105 -88
rect -40935 -190 -40795 190
rect -38715 88 -38695 4232
rect -38595 88 -38575 4232
rect -36405 4130 -36265 4320
rect -34185 4232 -34045 4320
rect -38715 -88 -38575 88
rect -43245 -4320 -43105 -4232
rect -40935 -4320 -40795 -4130
rect -38715 -4232 -38695 -88
rect -38595 -4232 -38575 -88
rect -36405 -190 -36265 190
rect -34185 88 -34165 4232
rect -34065 88 -34045 4232
rect -31875 4130 -31735 4320
rect -29655 4232 -29515 4320
rect -34185 -88 -34045 88
rect -38715 -4320 -38575 -4232
rect -36405 -4320 -36265 -4130
rect -34185 -4232 -34165 -88
rect -34065 -4232 -34045 -88
rect -31875 -190 -31735 190
rect -29655 88 -29635 4232
rect -29535 88 -29515 4232
rect -27345 4130 -27205 4320
rect -25125 4232 -24985 4320
rect -29655 -88 -29515 88
rect -34185 -4320 -34045 -4232
rect -31875 -4320 -31735 -4130
rect -29655 -4232 -29635 -88
rect -29535 -4232 -29515 -88
rect -27345 -190 -27205 190
rect -25125 88 -25105 4232
rect -25005 88 -24985 4232
rect -22815 4130 -22675 4320
rect -20595 4232 -20455 4320
rect -25125 -88 -24985 88
rect -29655 -4320 -29515 -4232
rect -27345 -4320 -27205 -4130
rect -25125 -4232 -25105 -88
rect -25005 -4232 -24985 -88
rect -22815 -190 -22675 190
rect -20595 88 -20575 4232
rect -20475 88 -20455 4232
rect -18285 4130 -18145 4320
rect -16065 4232 -15925 4320
rect -20595 -88 -20455 88
rect -25125 -4320 -24985 -4232
rect -22815 -4320 -22675 -4130
rect -20595 -4232 -20575 -88
rect -20475 -4232 -20455 -88
rect -18285 -190 -18145 190
rect -16065 88 -16045 4232
rect -15945 88 -15925 4232
rect -13755 4130 -13615 4320
rect -11535 4232 -11395 4320
rect -16065 -88 -15925 88
rect -20595 -4320 -20455 -4232
rect -18285 -4320 -18145 -4130
rect -16065 -4232 -16045 -88
rect -15945 -4232 -15925 -88
rect -13755 -190 -13615 190
rect -11535 88 -11515 4232
rect -11415 88 -11395 4232
rect -9225 4130 -9085 4320
rect -7005 4232 -6865 4320
rect -11535 -88 -11395 88
rect -16065 -4320 -15925 -4232
rect -13755 -4320 -13615 -4130
rect -11535 -4232 -11515 -88
rect -11415 -4232 -11395 -88
rect -9225 -190 -9085 190
rect -7005 88 -6985 4232
rect -6885 88 -6865 4232
rect -4695 4130 -4555 4320
rect -2475 4232 -2335 4320
rect -7005 -88 -6865 88
rect -11535 -4320 -11395 -4232
rect -9225 -4320 -9085 -4130
rect -7005 -4232 -6985 -88
rect -6885 -4232 -6865 -88
rect -4695 -190 -4555 190
rect -2475 88 -2455 4232
rect -2355 88 -2335 4232
rect -165 4130 -25 4320
rect 2055 4232 2195 4320
rect -2475 -88 -2335 88
rect -7005 -4320 -6865 -4232
rect -4695 -4320 -4555 -4130
rect -2475 -4232 -2455 -88
rect -2355 -4232 -2335 -88
rect -165 -190 -25 190
rect 2055 88 2075 4232
rect 2175 88 2195 4232
rect 4365 4130 4505 4320
rect 6585 4232 6725 4320
rect 2055 -88 2195 88
rect -2475 -4320 -2335 -4232
rect -165 -4320 -25 -4130
rect 2055 -4232 2075 -88
rect 2175 -4232 2195 -88
rect 4365 -190 4505 190
rect 6585 88 6605 4232
rect 6705 88 6725 4232
rect 8895 4130 9035 4320
rect 11115 4232 11255 4320
rect 6585 -88 6725 88
rect 2055 -4320 2195 -4232
rect 4365 -4320 4505 -4130
rect 6585 -4232 6605 -88
rect 6705 -4232 6725 -88
rect 8895 -190 9035 190
rect 11115 88 11135 4232
rect 11235 88 11255 4232
rect 13425 4130 13565 4320
rect 15645 4232 15785 4320
rect 11115 -88 11255 88
rect 6585 -4320 6725 -4232
rect 8895 -4320 9035 -4130
rect 11115 -4232 11135 -88
rect 11235 -4232 11255 -88
rect 13425 -190 13565 190
rect 15645 88 15665 4232
rect 15765 88 15785 4232
rect 17955 4130 18095 4320
rect 20175 4232 20315 4320
rect 15645 -88 15785 88
rect 11115 -4320 11255 -4232
rect 13425 -4320 13565 -4130
rect 15645 -4232 15665 -88
rect 15765 -4232 15785 -88
rect 17955 -190 18095 190
rect 20175 88 20195 4232
rect 20295 88 20315 4232
rect 22485 4130 22625 4320
rect 24705 4232 24845 4320
rect 20175 -88 20315 88
rect 15645 -4320 15785 -4232
rect 17955 -4320 18095 -4130
rect 20175 -4232 20195 -88
rect 20295 -4232 20315 -88
rect 22485 -190 22625 190
rect 24705 88 24725 4232
rect 24825 88 24845 4232
rect 27015 4130 27155 4320
rect 29235 4232 29375 4320
rect 24705 -88 24845 88
rect 20175 -4320 20315 -4232
rect 22485 -4320 22625 -4130
rect 24705 -4232 24725 -88
rect 24825 -4232 24845 -88
rect 27015 -190 27155 190
rect 29235 88 29255 4232
rect 29355 88 29375 4232
rect 31545 4130 31685 4320
rect 33765 4232 33905 4320
rect 29235 -88 29375 88
rect 24705 -4320 24845 -4232
rect 27015 -4320 27155 -4130
rect 29235 -4232 29255 -88
rect 29355 -4232 29375 -88
rect 31545 -190 31685 190
rect 33765 88 33785 4232
rect 33885 88 33905 4232
rect 36075 4130 36215 4320
rect 38295 4232 38435 4320
rect 33765 -88 33905 88
rect 29235 -4320 29375 -4232
rect 31545 -4320 31685 -4130
rect 33765 -4232 33785 -88
rect 33885 -4232 33905 -88
rect 36075 -190 36215 190
rect 38295 88 38315 4232
rect 38415 88 38435 4232
rect 40605 4130 40745 4320
rect 42825 4232 42965 4320
rect 38295 -88 38435 88
rect 33765 -4320 33905 -4232
rect 36075 -4320 36215 -4130
rect 38295 -4232 38315 -88
rect 38415 -4232 38435 -88
rect 40605 -190 40745 190
rect 42825 88 42845 4232
rect 42945 88 42965 4232
rect 45135 4130 45275 4320
rect 47355 4232 47495 4320
rect 42825 -88 42965 88
rect 38295 -4320 38435 -4232
rect 40605 -4320 40745 -4130
rect 42825 -4232 42845 -88
rect 42945 -4232 42965 -88
rect 45135 -190 45275 190
rect 47355 88 47375 4232
rect 47475 88 47495 4232
rect 49665 4130 49805 4320
rect 51885 4232 52025 4320
rect 47355 -88 47495 88
rect 42825 -4320 42965 -4232
rect 45135 -4320 45275 -4130
rect 47355 -4232 47375 -88
rect 47475 -4232 47495 -88
rect 49665 -190 49805 190
rect 51885 88 51905 4232
rect 52005 88 52025 4232
rect 54195 4130 54335 4320
rect 56415 4232 56555 4320
rect 51885 -88 52025 88
rect 47355 -4320 47495 -4232
rect 49665 -4320 49805 -4130
rect 51885 -4232 51905 -88
rect 52005 -4232 52025 -88
rect 54195 -190 54335 190
rect 56415 88 56435 4232
rect 56535 88 56555 4232
rect 58725 4130 58865 4320
rect 60945 4232 61085 4320
rect 56415 -88 56555 88
rect 51885 -4320 52025 -4232
rect 54195 -4320 54335 -4130
rect 56415 -4232 56435 -88
rect 56535 -4232 56555 -88
rect 58725 -190 58865 190
rect 60945 88 60965 4232
rect 61065 88 61085 4232
rect 63255 4130 63395 4320
rect 65475 4232 65615 4320
rect 60945 -88 61085 88
rect 56415 -4320 56555 -4232
rect 58725 -4320 58865 -4130
rect 60945 -4232 60965 -88
rect 61065 -4232 61085 -88
rect 63255 -190 63395 190
rect 65475 88 65495 4232
rect 65595 88 65615 4232
rect 67785 4130 67925 4320
rect 70005 4232 70145 4320
rect 65475 -88 65615 88
rect 60945 -4320 61085 -4232
rect 63255 -4320 63395 -4130
rect 65475 -4232 65495 -88
rect 65595 -4232 65615 -88
rect 67785 -190 67925 190
rect 70005 88 70025 4232
rect 70125 88 70145 4232
rect 72315 4130 72455 4320
rect 74535 4232 74675 4320
rect 70005 -88 70145 88
rect 65475 -4320 65615 -4232
rect 67785 -4320 67925 -4130
rect 70005 -4232 70025 -88
rect 70125 -4232 70145 -88
rect 72315 -190 72455 190
rect 74535 88 74555 4232
rect 74655 88 74675 4232
rect 76845 4130 76985 4320
rect 79065 4232 79205 4320
rect 74535 -88 74675 88
rect 70005 -4320 70145 -4232
rect 72315 -4320 72455 -4130
rect 74535 -4232 74555 -88
rect 74655 -4232 74675 -88
rect 76845 -190 76985 190
rect 79065 88 79085 4232
rect 79185 88 79205 4232
rect 79065 -88 79205 88
rect 74535 -4320 74675 -4232
rect 76845 -4320 76985 -4130
rect 79065 -4232 79085 -88
rect 79185 -4232 79205 -88
rect 79065 -4320 79205 -4232
<< properties >>
string parameters w 20.00 l 20.00 val 413.6 carea 1.00 cperi 0.17 nx 35 ny 2 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
