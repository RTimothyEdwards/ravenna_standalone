magic
tech EFXH018D
magscale 1 2
timestamp 1565723183
<< mimcap >>
rect -124405 6290 -120405 6320
rect -124405 2350 -124375 6290
rect -120435 2350 -120405 6290
rect -124405 2320 -120405 2350
rect -119875 6290 -115875 6320
rect -119875 2350 -119845 6290
rect -115905 2350 -115875 6290
rect -119875 2320 -115875 2350
rect -115345 6290 -111345 6320
rect -115345 2350 -115315 6290
rect -111375 2350 -111345 6290
rect -115345 2320 -111345 2350
rect -110815 6290 -106815 6320
rect -110815 2350 -110785 6290
rect -106845 2350 -106815 6290
rect -110815 2320 -106815 2350
rect -106285 6290 -102285 6320
rect -106285 2350 -106255 6290
rect -102315 2350 -102285 6290
rect -106285 2320 -102285 2350
rect -101755 6290 -97755 6320
rect -101755 2350 -101725 6290
rect -97785 2350 -97755 6290
rect -101755 2320 -97755 2350
rect -97225 6290 -93225 6320
rect -97225 2350 -97195 6290
rect -93255 2350 -93225 6290
rect -97225 2320 -93225 2350
rect -92695 6290 -88695 6320
rect -92695 2350 -92665 6290
rect -88725 2350 -88695 6290
rect -92695 2320 -88695 2350
rect -88165 6290 -84165 6320
rect -88165 2350 -88135 6290
rect -84195 2350 -84165 6290
rect -88165 2320 -84165 2350
rect -83635 6290 -79635 6320
rect -83635 2350 -83605 6290
rect -79665 2350 -79635 6290
rect -83635 2320 -79635 2350
rect -79105 6290 -75105 6320
rect -79105 2350 -79075 6290
rect -75135 2350 -75105 6290
rect -79105 2320 -75105 2350
rect -74575 6290 -70575 6320
rect -74575 2350 -74545 6290
rect -70605 2350 -70575 6290
rect -74575 2320 -70575 2350
rect -70045 6290 -66045 6320
rect -70045 2350 -70015 6290
rect -66075 2350 -66045 6290
rect -70045 2320 -66045 2350
rect -65515 6290 -61515 6320
rect -65515 2350 -65485 6290
rect -61545 2350 -61515 6290
rect -65515 2320 -61515 2350
rect -60985 6290 -56985 6320
rect -60985 2350 -60955 6290
rect -57015 2350 -56985 6290
rect -60985 2320 -56985 2350
rect -56455 6290 -52455 6320
rect -56455 2350 -56425 6290
rect -52485 2350 -52455 6290
rect -56455 2320 -52455 2350
rect -51925 6290 -47925 6320
rect -51925 2350 -51895 6290
rect -47955 2350 -47925 6290
rect -51925 2320 -47925 2350
rect -47395 6290 -43395 6320
rect -47395 2350 -47365 6290
rect -43425 2350 -43395 6290
rect -47395 2320 -43395 2350
rect -42865 6290 -38865 6320
rect -42865 2350 -42835 6290
rect -38895 2350 -38865 6290
rect -42865 2320 -38865 2350
rect -38335 6290 -34335 6320
rect -38335 2350 -38305 6290
rect -34365 2350 -34335 6290
rect -38335 2320 -34335 2350
rect -33805 6290 -29805 6320
rect -33805 2350 -33775 6290
rect -29835 2350 -29805 6290
rect -33805 2320 -29805 2350
rect -29275 6290 -25275 6320
rect -29275 2350 -29245 6290
rect -25305 2350 -25275 6290
rect -29275 2320 -25275 2350
rect -24745 6290 -20745 6320
rect -24745 2350 -24715 6290
rect -20775 2350 -20745 6290
rect -24745 2320 -20745 2350
rect -20215 6290 -16215 6320
rect -20215 2350 -20185 6290
rect -16245 2350 -16215 6290
rect -20215 2320 -16215 2350
rect -15685 6290 -11685 6320
rect -15685 2350 -15655 6290
rect -11715 2350 -11685 6290
rect -15685 2320 -11685 2350
rect -11155 6290 -7155 6320
rect -11155 2350 -11125 6290
rect -7185 2350 -7155 6290
rect -11155 2320 -7155 2350
rect -6625 6290 -2625 6320
rect -6625 2350 -6595 6290
rect -2655 2350 -2625 6290
rect -6625 2320 -2625 2350
rect -2095 6290 1905 6320
rect -2095 2350 -2065 6290
rect 1875 2350 1905 6290
rect -2095 2320 1905 2350
rect 2435 6290 6435 6320
rect 2435 2350 2465 6290
rect 6405 2350 6435 6290
rect 2435 2320 6435 2350
rect 6965 6290 10965 6320
rect 6965 2350 6995 6290
rect 10935 2350 10965 6290
rect 6965 2320 10965 2350
rect 11495 6290 15495 6320
rect 11495 2350 11525 6290
rect 15465 2350 15495 6290
rect 11495 2320 15495 2350
rect 16025 6290 20025 6320
rect 16025 2350 16055 6290
rect 19995 2350 20025 6290
rect 16025 2320 20025 2350
rect 20555 6290 24555 6320
rect 20555 2350 20585 6290
rect 24525 2350 24555 6290
rect 20555 2320 24555 2350
rect 25085 6290 29085 6320
rect 25085 2350 25115 6290
rect 29055 2350 29085 6290
rect 25085 2320 29085 2350
rect 29615 6290 33615 6320
rect 29615 2350 29645 6290
rect 33585 2350 33615 6290
rect 29615 2320 33615 2350
rect 34145 6290 38145 6320
rect 34145 2350 34175 6290
rect 38115 2350 38145 6290
rect 34145 2320 38145 2350
rect 38675 6290 42675 6320
rect 38675 2350 38705 6290
rect 42645 2350 42675 6290
rect 38675 2320 42675 2350
rect 43205 6290 47205 6320
rect 43205 2350 43235 6290
rect 47175 2350 47205 6290
rect 43205 2320 47205 2350
rect 47735 6290 51735 6320
rect 47735 2350 47765 6290
rect 51705 2350 51735 6290
rect 47735 2320 51735 2350
rect 52265 6290 56265 6320
rect 52265 2350 52295 6290
rect 56235 2350 56265 6290
rect 52265 2320 56265 2350
rect 56795 6290 60795 6320
rect 56795 2350 56825 6290
rect 60765 2350 60795 6290
rect 56795 2320 60795 2350
rect 61325 6290 65325 6320
rect 61325 2350 61355 6290
rect 65295 2350 65325 6290
rect 61325 2320 65325 2350
rect 65855 6290 69855 6320
rect 65855 2350 65885 6290
rect 69825 2350 69855 6290
rect 65855 2320 69855 2350
rect 70385 6290 74385 6320
rect 70385 2350 70415 6290
rect 74355 2350 74385 6290
rect 70385 2320 74385 2350
rect 74915 6290 78915 6320
rect 74915 2350 74945 6290
rect 78885 2350 78915 6290
rect 74915 2320 78915 2350
rect 79445 6290 83445 6320
rect 79445 2350 79475 6290
rect 83415 2350 83445 6290
rect 79445 2320 83445 2350
rect 83975 6290 87975 6320
rect 83975 2350 84005 6290
rect 87945 2350 87975 6290
rect 83975 2320 87975 2350
rect 88505 6290 92505 6320
rect 88505 2350 88535 6290
rect 92475 2350 92505 6290
rect 88505 2320 92505 2350
rect 93035 6290 97035 6320
rect 93035 2350 93065 6290
rect 97005 2350 97035 6290
rect 93035 2320 97035 2350
rect 97565 6290 101565 6320
rect 97565 2350 97595 6290
rect 101535 2350 101565 6290
rect 97565 2320 101565 2350
rect 102095 6290 106095 6320
rect 102095 2350 102125 6290
rect 106065 2350 106095 6290
rect 102095 2320 106095 2350
rect 106625 6290 110625 6320
rect 106625 2350 106655 6290
rect 110595 2350 110625 6290
rect 106625 2320 110625 2350
rect 111155 6290 115155 6320
rect 111155 2350 111185 6290
rect 115125 2350 115155 6290
rect 111155 2320 115155 2350
rect 115685 6290 119685 6320
rect 115685 2350 115715 6290
rect 119655 2350 119685 6290
rect 115685 2320 119685 2350
rect 120215 6290 124215 6320
rect 120215 2350 120245 6290
rect 124185 2350 124215 6290
rect 120215 2320 124215 2350
rect -124405 1970 -120405 2000
rect -124405 -1970 -124375 1970
rect -120435 -1970 -120405 1970
rect -124405 -2000 -120405 -1970
rect -119875 1970 -115875 2000
rect -119875 -1970 -119845 1970
rect -115905 -1970 -115875 1970
rect -119875 -2000 -115875 -1970
rect -115345 1970 -111345 2000
rect -115345 -1970 -115315 1970
rect -111375 -1970 -111345 1970
rect -115345 -2000 -111345 -1970
rect -110815 1970 -106815 2000
rect -110815 -1970 -110785 1970
rect -106845 -1970 -106815 1970
rect -110815 -2000 -106815 -1970
rect -106285 1970 -102285 2000
rect -106285 -1970 -106255 1970
rect -102315 -1970 -102285 1970
rect -106285 -2000 -102285 -1970
rect -101755 1970 -97755 2000
rect -101755 -1970 -101725 1970
rect -97785 -1970 -97755 1970
rect -101755 -2000 -97755 -1970
rect -97225 1970 -93225 2000
rect -97225 -1970 -97195 1970
rect -93255 -1970 -93225 1970
rect -97225 -2000 -93225 -1970
rect -92695 1970 -88695 2000
rect -92695 -1970 -92665 1970
rect -88725 -1970 -88695 1970
rect -92695 -2000 -88695 -1970
rect -88165 1970 -84165 2000
rect -88165 -1970 -88135 1970
rect -84195 -1970 -84165 1970
rect -88165 -2000 -84165 -1970
rect -83635 1970 -79635 2000
rect -83635 -1970 -83605 1970
rect -79665 -1970 -79635 1970
rect -83635 -2000 -79635 -1970
rect -79105 1970 -75105 2000
rect -79105 -1970 -79075 1970
rect -75135 -1970 -75105 1970
rect -79105 -2000 -75105 -1970
rect -74575 1970 -70575 2000
rect -74575 -1970 -74545 1970
rect -70605 -1970 -70575 1970
rect -74575 -2000 -70575 -1970
rect -70045 1970 -66045 2000
rect -70045 -1970 -70015 1970
rect -66075 -1970 -66045 1970
rect -70045 -2000 -66045 -1970
rect -65515 1970 -61515 2000
rect -65515 -1970 -65485 1970
rect -61545 -1970 -61515 1970
rect -65515 -2000 -61515 -1970
rect -60985 1970 -56985 2000
rect -60985 -1970 -60955 1970
rect -57015 -1970 -56985 1970
rect -60985 -2000 -56985 -1970
rect -56455 1970 -52455 2000
rect -56455 -1970 -56425 1970
rect -52485 -1970 -52455 1970
rect -56455 -2000 -52455 -1970
rect -51925 1970 -47925 2000
rect -51925 -1970 -51895 1970
rect -47955 -1970 -47925 1970
rect -51925 -2000 -47925 -1970
rect -47395 1970 -43395 2000
rect -47395 -1970 -47365 1970
rect -43425 -1970 -43395 1970
rect -47395 -2000 -43395 -1970
rect -42865 1970 -38865 2000
rect -42865 -1970 -42835 1970
rect -38895 -1970 -38865 1970
rect -42865 -2000 -38865 -1970
rect -38335 1970 -34335 2000
rect -38335 -1970 -38305 1970
rect -34365 -1970 -34335 1970
rect -38335 -2000 -34335 -1970
rect -33805 1970 -29805 2000
rect -33805 -1970 -33775 1970
rect -29835 -1970 -29805 1970
rect -33805 -2000 -29805 -1970
rect -29275 1970 -25275 2000
rect -29275 -1970 -29245 1970
rect -25305 -1970 -25275 1970
rect -29275 -2000 -25275 -1970
rect -24745 1970 -20745 2000
rect -24745 -1970 -24715 1970
rect -20775 -1970 -20745 1970
rect -24745 -2000 -20745 -1970
rect -20215 1970 -16215 2000
rect -20215 -1970 -20185 1970
rect -16245 -1970 -16215 1970
rect -20215 -2000 -16215 -1970
rect -15685 1970 -11685 2000
rect -15685 -1970 -15655 1970
rect -11715 -1970 -11685 1970
rect -15685 -2000 -11685 -1970
rect -11155 1970 -7155 2000
rect -11155 -1970 -11125 1970
rect -7185 -1970 -7155 1970
rect -11155 -2000 -7155 -1970
rect -6625 1970 -2625 2000
rect -6625 -1970 -6595 1970
rect -2655 -1970 -2625 1970
rect -6625 -2000 -2625 -1970
rect -2095 1970 1905 2000
rect -2095 -1970 -2065 1970
rect 1875 -1970 1905 1970
rect -2095 -2000 1905 -1970
rect 2435 1970 6435 2000
rect 2435 -1970 2465 1970
rect 6405 -1970 6435 1970
rect 2435 -2000 6435 -1970
rect 6965 1970 10965 2000
rect 6965 -1970 6995 1970
rect 10935 -1970 10965 1970
rect 6965 -2000 10965 -1970
rect 11495 1970 15495 2000
rect 11495 -1970 11525 1970
rect 15465 -1970 15495 1970
rect 11495 -2000 15495 -1970
rect 16025 1970 20025 2000
rect 16025 -1970 16055 1970
rect 19995 -1970 20025 1970
rect 16025 -2000 20025 -1970
rect 20555 1970 24555 2000
rect 20555 -1970 20585 1970
rect 24525 -1970 24555 1970
rect 20555 -2000 24555 -1970
rect 25085 1970 29085 2000
rect 25085 -1970 25115 1970
rect 29055 -1970 29085 1970
rect 25085 -2000 29085 -1970
rect 29615 1970 33615 2000
rect 29615 -1970 29645 1970
rect 33585 -1970 33615 1970
rect 29615 -2000 33615 -1970
rect 34145 1970 38145 2000
rect 34145 -1970 34175 1970
rect 38115 -1970 38145 1970
rect 34145 -2000 38145 -1970
rect 38675 1970 42675 2000
rect 38675 -1970 38705 1970
rect 42645 -1970 42675 1970
rect 38675 -2000 42675 -1970
rect 43205 1970 47205 2000
rect 43205 -1970 43235 1970
rect 47175 -1970 47205 1970
rect 43205 -2000 47205 -1970
rect 47735 1970 51735 2000
rect 47735 -1970 47765 1970
rect 51705 -1970 51735 1970
rect 47735 -2000 51735 -1970
rect 52265 1970 56265 2000
rect 52265 -1970 52295 1970
rect 56235 -1970 56265 1970
rect 52265 -2000 56265 -1970
rect 56795 1970 60795 2000
rect 56795 -1970 56825 1970
rect 60765 -1970 60795 1970
rect 56795 -2000 60795 -1970
rect 61325 1970 65325 2000
rect 61325 -1970 61355 1970
rect 65295 -1970 65325 1970
rect 61325 -2000 65325 -1970
rect 65855 1970 69855 2000
rect 65855 -1970 65885 1970
rect 69825 -1970 69855 1970
rect 65855 -2000 69855 -1970
rect 70385 1970 74385 2000
rect 70385 -1970 70415 1970
rect 74355 -1970 74385 1970
rect 70385 -2000 74385 -1970
rect 74915 1970 78915 2000
rect 74915 -1970 74945 1970
rect 78885 -1970 78915 1970
rect 74915 -2000 78915 -1970
rect 79445 1970 83445 2000
rect 79445 -1970 79475 1970
rect 83415 -1970 83445 1970
rect 79445 -2000 83445 -1970
rect 83975 1970 87975 2000
rect 83975 -1970 84005 1970
rect 87945 -1970 87975 1970
rect 83975 -2000 87975 -1970
rect 88505 1970 92505 2000
rect 88505 -1970 88535 1970
rect 92475 -1970 92505 1970
rect 88505 -2000 92505 -1970
rect 93035 1970 97035 2000
rect 93035 -1970 93065 1970
rect 97005 -1970 97035 1970
rect 93035 -2000 97035 -1970
rect 97565 1970 101565 2000
rect 97565 -1970 97595 1970
rect 101535 -1970 101565 1970
rect 97565 -2000 101565 -1970
rect 102095 1970 106095 2000
rect 102095 -1970 102125 1970
rect 106065 -1970 106095 1970
rect 102095 -2000 106095 -1970
rect 106625 1970 110625 2000
rect 106625 -1970 106655 1970
rect 110595 -1970 110625 1970
rect 106625 -2000 110625 -1970
rect 111155 1970 115155 2000
rect 111155 -1970 111185 1970
rect 115125 -1970 115155 1970
rect 111155 -2000 115155 -1970
rect 115685 1970 119685 2000
rect 115685 -1970 115715 1970
rect 119655 -1970 119685 1970
rect 115685 -2000 119685 -1970
rect 120215 1970 124215 2000
rect 120215 -1970 120245 1970
rect 124185 -1970 124215 1970
rect 120215 -2000 124215 -1970
rect -124405 -2350 -120405 -2320
rect -124405 -6290 -124375 -2350
rect -120435 -6290 -120405 -2350
rect -124405 -6320 -120405 -6290
rect -119875 -2350 -115875 -2320
rect -119875 -6290 -119845 -2350
rect -115905 -6290 -115875 -2350
rect -119875 -6320 -115875 -6290
rect -115345 -2350 -111345 -2320
rect -115345 -6290 -115315 -2350
rect -111375 -6290 -111345 -2350
rect -115345 -6320 -111345 -6290
rect -110815 -2350 -106815 -2320
rect -110815 -6290 -110785 -2350
rect -106845 -6290 -106815 -2350
rect -110815 -6320 -106815 -6290
rect -106285 -2350 -102285 -2320
rect -106285 -6290 -106255 -2350
rect -102315 -6290 -102285 -2350
rect -106285 -6320 -102285 -6290
rect -101755 -2350 -97755 -2320
rect -101755 -6290 -101725 -2350
rect -97785 -6290 -97755 -2350
rect -101755 -6320 -97755 -6290
rect -97225 -2350 -93225 -2320
rect -97225 -6290 -97195 -2350
rect -93255 -6290 -93225 -2350
rect -97225 -6320 -93225 -6290
rect -92695 -2350 -88695 -2320
rect -92695 -6290 -92665 -2350
rect -88725 -6290 -88695 -2350
rect -92695 -6320 -88695 -6290
rect -88165 -2350 -84165 -2320
rect -88165 -6290 -88135 -2350
rect -84195 -6290 -84165 -2350
rect -88165 -6320 -84165 -6290
rect -83635 -2350 -79635 -2320
rect -83635 -6290 -83605 -2350
rect -79665 -6290 -79635 -2350
rect -83635 -6320 -79635 -6290
rect -79105 -2350 -75105 -2320
rect -79105 -6290 -79075 -2350
rect -75135 -6290 -75105 -2350
rect -79105 -6320 -75105 -6290
rect -74575 -2350 -70575 -2320
rect -74575 -6290 -74545 -2350
rect -70605 -6290 -70575 -2350
rect -74575 -6320 -70575 -6290
rect -70045 -2350 -66045 -2320
rect -70045 -6290 -70015 -2350
rect -66075 -6290 -66045 -2350
rect -70045 -6320 -66045 -6290
rect -65515 -2350 -61515 -2320
rect -65515 -6290 -65485 -2350
rect -61545 -6290 -61515 -2350
rect -65515 -6320 -61515 -6290
rect -60985 -2350 -56985 -2320
rect -60985 -6290 -60955 -2350
rect -57015 -6290 -56985 -2350
rect -60985 -6320 -56985 -6290
rect -56455 -2350 -52455 -2320
rect -56455 -6290 -56425 -2350
rect -52485 -6290 -52455 -2350
rect -56455 -6320 -52455 -6290
rect -51925 -2350 -47925 -2320
rect -51925 -6290 -51895 -2350
rect -47955 -6290 -47925 -2350
rect -51925 -6320 -47925 -6290
rect -47395 -2350 -43395 -2320
rect -47395 -6290 -47365 -2350
rect -43425 -6290 -43395 -2350
rect -47395 -6320 -43395 -6290
rect -42865 -2350 -38865 -2320
rect -42865 -6290 -42835 -2350
rect -38895 -6290 -38865 -2350
rect -42865 -6320 -38865 -6290
rect -38335 -2350 -34335 -2320
rect -38335 -6290 -38305 -2350
rect -34365 -6290 -34335 -2350
rect -38335 -6320 -34335 -6290
rect -33805 -2350 -29805 -2320
rect -33805 -6290 -33775 -2350
rect -29835 -6290 -29805 -2350
rect -33805 -6320 -29805 -6290
rect -29275 -2350 -25275 -2320
rect -29275 -6290 -29245 -2350
rect -25305 -6290 -25275 -2350
rect -29275 -6320 -25275 -6290
rect -24745 -2350 -20745 -2320
rect -24745 -6290 -24715 -2350
rect -20775 -6290 -20745 -2350
rect -24745 -6320 -20745 -6290
rect -20215 -2350 -16215 -2320
rect -20215 -6290 -20185 -2350
rect -16245 -6290 -16215 -2350
rect -20215 -6320 -16215 -6290
rect -15685 -2350 -11685 -2320
rect -15685 -6290 -15655 -2350
rect -11715 -6290 -11685 -2350
rect -15685 -6320 -11685 -6290
rect -11155 -2350 -7155 -2320
rect -11155 -6290 -11125 -2350
rect -7185 -6290 -7155 -2350
rect -11155 -6320 -7155 -6290
rect -6625 -2350 -2625 -2320
rect -6625 -6290 -6595 -2350
rect -2655 -6290 -2625 -2350
rect -6625 -6320 -2625 -6290
rect -2095 -2350 1905 -2320
rect -2095 -6290 -2065 -2350
rect 1875 -6290 1905 -2350
rect -2095 -6320 1905 -6290
rect 2435 -2350 6435 -2320
rect 2435 -6290 2465 -2350
rect 6405 -6290 6435 -2350
rect 2435 -6320 6435 -6290
rect 6965 -2350 10965 -2320
rect 6965 -6290 6995 -2350
rect 10935 -6290 10965 -2350
rect 6965 -6320 10965 -6290
rect 11495 -2350 15495 -2320
rect 11495 -6290 11525 -2350
rect 15465 -6290 15495 -2350
rect 11495 -6320 15495 -6290
rect 16025 -2350 20025 -2320
rect 16025 -6290 16055 -2350
rect 19995 -6290 20025 -2350
rect 16025 -6320 20025 -6290
rect 20555 -2350 24555 -2320
rect 20555 -6290 20585 -2350
rect 24525 -6290 24555 -2350
rect 20555 -6320 24555 -6290
rect 25085 -2350 29085 -2320
rect 25085 -6290 25115 -2350
rect 29055 -6290 29085 -2350
rect 25085 -6320 29085 -6290
rect 29615 -2350 33615 -2320
rect 29615 -6290 29645 -2350
rect 33585 -6290 33615 -2350
rect 29615 -6320 33615 -6290
rect 34145 -2350 38145 -2320
rect 34145 -6290 34175 -2350
rect 38115 -6290 38145 -2350
rect 34145 -6320 38145 -6290
rect 38675 -2350 42675 -2320
rect 38675 -6290 38705 -2350
rect 42645 -6290 42675 -2350
rect 38675 -6320 42675 -6290
rect 43205 -2350 47205 -2320
rect 43205 -6290 43235 -2350
rect 47175 -6290 47205 -2350
rect 43205 -6320 47205 -6290
rect 47735 -2350 51735 -2320
rect 47735 -6290 47765 -2350
rect 51705 -6290 51735 -2350
rect 47735 -6320 51735 -6290
rect 52265 -2350 56265 -2320
rect 52265 -6290 52295 -2350
rect 56235 -6290 56265 -2350
rect 52265 -6320 56265 -6290
rect 56795 -2350 60795 -2320
rect 56795 -6290 56825 -2350
rect 60765 -6290 60795 -2350
rect 56795 -6320 60795 -6290
rect 61325 -2350 65325 -2320
rect 61325 -6290 61355 -2350
rect 65295 -6290 65325 -2350
rect 61325 -6320 65325 -6290
rect 65855 -2350 69855 -2320
rect 65855 -6290 65885 -2350
rect 69825 -6290 69855 -2350
rect 65855 -6320 69855 -6290
rect 70385 -2350 74385 -2320
rect 70385 -6290 70415 -2350
rect 74355 -6290 74385 -2350
rect 70385 -6320 74385 -6290
rect 74915 -2350 78915 -2320
rect 74915 -6290 74945 -2350
rect 78885 -6290 78915 -2350
rect 74915 -6320 78915 -6290
rect 79445 -2350 83445 -2320
rect 79445 -6290 79475 -2350
rect 83415 -6290 83445 -2350
rect 79445 -6320 83445 -6290
rect 83975 -2350 87975 -2320
rect 83975 -6290 84005 -2350
rect 87945 -6290 87975 -2350
rect 83975 -6320 87975 -6290
rect 88505 -2350 92505 -2320
rect 88505 -6290 88535 -2350
rect 92475 -6290 92505 -2350
rect 88505 -6320 92505 -6290
rect 93035 -2350 97035 -2320
rect 93035 -6290 93065 -2350
rect 97005 -6290 97035 -2350
rect 93035 -6320 97035 -6290
rect 97565 -2350 101565 -2320
rect 97565 -6290 97595 -2350
rect 101535 -6290 101565 -2350
rect 97565 -6320 101565 -6290
rect 102095 -2350 106095 -2320
rect 102095 -6290 102125 -2350
rect 106065 -6290 106095 -2350
rect 102095 -6320 106095 -6290
rect 106625 -2350 110625 -2320
rect 106625 -6290 106655 -2350
rect 110595 -6290 110625 -2350
rect 106625 -6320 110625 -6290
rect 111155 -2350 115155 -2320
rect 111155 -6290 111185 -2350
rect 115125 -6290 115155 -2350
rect 111155 -6320 115155 -6290
rect 115685 -2350 119685 -2320
rect 115685 -6290 115715 -2350
rect 119655 -6290 119685 -2350
rect 115685 -6320 119685 -6290
rect 120215 -2350 124215 -2320
rect 120215 -6290 120245 -2350
rect 124185 -6290 124215 -2350
rect 120215 -6320 124215 -6290
<< mimcapcontact >>
rect -124375 2350 -120435 6290
rect -119845 2350 -115905 6290
rect -115315 2350 -111375 6290
rect -110785 2350 -106845 6290
rect -106255 2350 -102315 6290
rect -101725 2350 -97785 6290
rect -97195 2350 -93255 6290
rect -92665 2350 -88725 6290
rect -88135 2350 -84195 6290
rect -83605 2350 -79665 6290
rect -79075 2350 -75135 6290
rect -74545 2350 -70605 6290
rect -70015 2350 -66075 6290
rect -65485 2350 -61545 6290
rect -60955 2350 -57015 6290
rect -56425 2350 -52485 6290
rect -51895 2350 -47955 6290
rect -47365 2350 -43425 6290
rect -42835 2350 -38895 6290
rect -38305 2350 -34365 6290
rect -33775 2350 -29835 6290
rect -29245 2350 -25305 6290
rect -24715 2350 -20775 6290
rect -20185 2350 -16245 6290
rect -15655 2350 -11715 6290
rect -11125 2350 -7185 6290
rect -6595 2350 -2655 6290
rect -2065 2350 1875 6290
rect 2465 2350 6405 6290
rect 6995 2350 10935 6290
rect 11525 2350 15465 6290
rect 16055 2350 19995 6290
rect 20585 2350 24525 6290
rect 25115 2350 29055 6290
rect 29645 2350 33585 6290
rect 34175 2350 38115 6290
rect 38705 2350 42645 6290
rect 43235 2350 47175 6290
rect 47765 2350 51705 6290
rect 52295 2350 56235 6290
rect 56825 2350 60765 6290
rect 61355 2350 65295 6290
rect 65885 2350 69825 6290
rect 70415 2350 74355 6290
rect 74945 2350 78885 6290
rect 79475 2350 83415 6290
rect 84005 2350 87945 6290
rect 88535 2350 92475 6290
rect 93065 2350 97005 6290
rect 97595 2350 101535 6290
rect 102125 2350 106065 6290
rect 106655 2350 110595 6290
rect 111185 2350 115125 6290
rect 115715 2350 119655 6290
rect 120245 2350 124185 6290
rect -124375 -1970 -120435 1970
rect -119845 -1970 -115905 1970
rect -115315 -1970 -111375 1970
rect -110785 -1970 -106845 1970
rect -106255 -1970 -102315 1970
rect -101725 -1970 -97785 1970
rect -97195 -1970 -93255 1970
rect -92665 -1970 -88725 1970
rect -88135 -1970 -84195 1970
rect -83605 -1970 -79665 1970
rect -79075 -1970 -75135 1970
rect -74545 -1970 -70605 1970
rect -70015 -1970 -66075 1970
rect -65485 -1970 -61545 1970
rect -60955 -1970 -57015 1970
rect -56425 -1970 -52485 1970
rect -51895 -1970 -47955 1970
rect -47365 -1970 -43425 1970
rect -42835 -1970 -38895 1970
rect -38305 -1970 -34365 1970
rect -33775 -1970 -29835 1970
rect -29245 -1970 -25305 1970
rect -24715 -1970 -20775 1970
rect -20185 -1970 -16245 1970
rect -15655 -1970 -11715 1970
rect -11125 -1970 -7185 1970
rect -6595 -1970 -2655 1970
rect -2065 -1970 1875 1970
rect 2465 -1970 6405 1970
rect 6995 -1970 10935 1970
rect 11525 -1970 15465 1970
rect 16055 -1970 19995 1970
rect 20585 -1970 24525 1970
rect 25115 -1970 29055 1970
rect 29645 -1970 33585 1970
rect 34175 -1970 38115 1970
rect 38705 -1970 42645 1970
rect 43235 -1970 47175 1970
rect 47765 -1970 51705 1970
rect 52295 -1970 56235 1970
rect 56825 -1970 60765 1970
rect 61355 -1970 65295 1970
rect 65885 -1970 69825 1970
rect 70415 -1970 74355 1970
rect 74945 -1970 78885 1970
rect 79475 -1970 83415 1970
rect 84005 -1970 87945 1970
rect 88535 -1970 92475 1970
rect 93065 -1970 97005 1970
rect 97595 -1970 101535 1970
rect 102125 -1970 106065 1970
rect 106655 -1970 110595 1970
rect 111185 -1970 115125 1970
rect 115715 -1970 119655 1970
rect 120245 -1970 124185 1970
rect -124375 -6290 -120435 -2350
rect -119845 -6290 -115905 -2350
rect -115315 -6290 -111375 -2350
rect -110785 -6290 -106845 -2350
rect -106255 -6290 -102315 -2350
rect -101725 -6290 -97785 -2350
rect -97195 -6290 -93255 -2350
rect -92665 -6290 -88725 -2350
rect -88135 -6290 -84195 -2350
rect -83605 -6290 -79665 -2350
rect -79075 -6290 -75135 -2350
rect -74545 -6290 -70605 -2350
rect -70015 -6290 -66075 -2350
rect -65485 -6290 -61545 -2350
rect -60955 -6290 -57015 -2350
rect -56425 -6290 -52485 -2350
rect -51895 -6290 -47955 -2350
rect -47365 -6290 -43425 -2350
rect -42835 -6290 -38895 -2350
rect -38305 -6290 -34365 -2350
rect -33775 -6290 -29835 -2350
rect -29245 -6290 -25305 -2350
rect -24715 -6290 -20775 -2350
rect -20185 -6290 -16245 -2350
rect -15655 -6290 -11715 -2350
rect -11125 -6290 -7185 -2350
rect -6595 -6290 -2655 -2350
rect -2065 -6290 1875 -2350
rect 2465 -6290 6405 -2350
rect 6995 -6290 10935 -2350
rect 11525 -6290 15465 -2350
rect 16055 -6290 19995 -2350
rect 20585 -6290 24525 -2350
rect 25115 -6290 29055 -2350
rect 29645 -6290 33585 -2350
rect 34175 -6290 38115 -2350
rect 38705 -6290 42645 -2350
rect 43235 -6290 47175 -2350
rect 47765 -6290 51705 -2350
rect 52295 -6290 56235 -2350
rect 56825 -6290 60765 -2350
rect 61355 -6290 65295 -2350
rect 65885 -6290 69825 -2350
rect 70415 -6290 74355 -2350
rect 74945 -6290 78885 -2350
rect 79475 -6290 83415 -2350
rect 84005 -6290 87945 -2350
rect 88535 -6290 92475 -2350
rect 93065 -6290 97005 -2350
rect 97595 -6290 101535 -2350
rect 102125 -6290 106065 -2350
rect 106655 -6290 110595 -2350
rect 111185 -6290 115125 -2350
rect 115715 -6290 119655 -2350
rect 120245 -6290 124185 -2350
<< metal4 >>
rect -124505 6392 -120115 6420
rect -124505 6320 -120235 6392
rect -124505 2320 -124405 6320
rect -120405 2320 -120235 6320
rect -124505 2248 -120235 2320
rect -120135 2248 -120115 6392
rect -124505 2220 -120115 2248
rect -119975 6392 -115585 6420
rect -119975 6320 -115705 6392
rect -119975 2320 -119875 6320
rect -115875 2320 -115705 6320
rect -119975 2248 -115705 2320
rect -115605 2248 -115585 6392
rect -119975 2220 -115585 2248
rect -115445 6392 -111055 6420
rect -115445 6320 -111175 6392
rect -115445 2320 -115345 6320
rect -111345 2320 -111175 6320
rect -115445 2248 -111175 2320
rect -111075 2248 -111055 6392
rect -115445 2220 -111055 2248
rect -110915 6392 -106525 6420
rect -110915 6320 -106645 6392
rect -110915 2320 -110815 6320
rect -106815 2320 -106645 6320
rect -110915 2248 -106645 2320
rect -106545 2248 -106525 6392
rect -110915 2220 -106525 2248
rect -106385 6392 -101995 6420
rect -106385 6320 -102115 6392
rect -106385 2320 -106285 6320
rect -102285 2320 -102115 6320
rect -106385 2248 -102115 2320
rect -102015 2248 -101995 6392
rect -106385 2220 -101995 2248
rect -101855 6392 -97465 6420
rect -101855 6320 -97585 6392
rect -101855 2320 -101755 6320
rect -97755 2320 -97585 6320
rect -101855 2248 -97585 2320
rect -97485 2248 -97465 6392
rect -101855 2220 -97465 2248
rect -97325 6392 -92935 6420
rect -97325 6320 -93055 6392
rect -97325 2320 -97225 6320
rect -93225 2320 -93055 6320
rect -97325 2248 -93055 2320
rect -92955 2248 -92935 6392
rect -97325 2220 -92935 2248
rect -92795 6392 -88405 6420
rect -92795 6320 -88525 6392
rect -92795 2320 -92695 6320
rect -88695 2320 -88525 6320
rect -92795 2248 -88525 2320
rect -88425 2248 -88405 6392
rect -92795 2220 -88405 2248
rect -88265 6392 -83875 6420
rect -88265 6320 -83995 6392
rect -88265 2320 -88165 6320
rect -84165 2320 -83995 6320
rect -88265 2248 -83995 2320
rect -83895 2248 -83875 6392
rect -88265 2220 -83875 2248
rect -83735 6392 -79345 6420
rect -83735 6320 -79465 6392
rect -83735 2320 -83635 6320
rect -79635 2320 -79465 6320
rect -83735 2248 -79465 2320
rect -79365 2248 -79345 6392
rect -83735 2220 -79345 2248
rect -79205 6392 -74815 6420
rect -79205 6320 -74935 6392
rect -79205 2320 -79105 6320
rect -75105 2320 -74935 6320
rect -79205 2248 -74935 2320
rect -74835 2248 -74815 6392
rect -79205 2220 -74815 2248
rect -74675 6392 -70285 6420
rect -74675 6320 -70405 6392
rect -74675 2320 -74575 6320
rect -70575 2320 -70405 6320
rect -74675 2248 -70405 2320
rect -70305 2248 -70285 6392
rect -74675 2220 -70285 2248
rect -70145 6392 -65755 6420
rect -70145 6320 -65875 6392
rect -70145 2320 -70045 6320
rect -66045 2320 -65875 6320
rect -70145 2248 -65875 2320
rect -65775 2248 -65755 6392
rect -70145 2220 -65755 2248
rect -65615 6392 -61225 6420
rect -65615 6320 -61345 6392
rect -65615 2320 -65515 6320
rect -61515 2320 -61345 6320
rect -65615 2248 -61345 2320
rect -61245 2248 -61225 6392
rect -65615 2220 -61225 2248
rect -61085 6392 -56695 6420
rect -61085 6320 -56815 6392
rect -61085 2320 -60985 6320
rect -56985 2320 -56815 6320
rect -61085 2248 -56815 2320
rect -56715 2248 -56695 6392
rect -61085 2220 -56695 2248
rect -56555 6392 -52165 6420
rect -56555 6320 -52285 6392
rect -56555 2320 -56455 6320
rect -52455 2320 -52285 6320
rect -56555 2248 -52285 2320
rect -52185 2248 -52165 6392
rect -56555 2220 -52165 2248
rect -52025 6392 -47635 6420
rect -52025 6320 -47755 6392
rect -52025 2320 -51925 6320
rect -47925 2320 -47755 6320
rect -52025 2248 -47755 2320
rect -47655 2248 -47635 6392
rect -52025 2220 -47635 2248
rect -47495 6392 -43105 6420
rect -47495 6320 -43225 6392
rect -47495 2320 -47395 6320
rect -43395 2320 -43225 6320
rect -47495 2248 -43225 2320
rect -43125 2248 -43105 6392
rect -47495 2220 -43105 2248
rect -42965 6392 -38575 6420
rect -42965 6320 -38695 6392
rect -42965 2320 -42865 6320
rect -38865 2320 -38695 6320
rect -42965 2248 -38695 2320
rect -38595 2248 -38575 6392
rect -42965 2220 -38575 2248
rect -38435 6392 -34045 6420
rect -38435 6320 -34165 6392
rect -38435 2320 -38335 6320
rect -34335 2320 -34165 6320
rect -38435 2248 -34165 2320
rect -34065 2248 -34045 6392
rect -38435 2220 -34045 2248
rect -33905 6392 -29515 6420
rect -33905 6320 -29635 6392
rect -33905 2320 -33805 6320
rect -29805 2320 -29635 6320
rect -33905 2248 -29635 2320
rect -29535 2248 -29515 6392
rect -33905 2220 -29515 2248
rect -29375 6392 -24985 6420
rect -29375 6320 -25105 6392
rect -29375 2320 -29275 6320
rect -25275 2320 -25105 6320
rect -29375 2248 -25105 2320
rect -25005 2248 -24985 6392
rect -29375 2220 -24985 2248
rect -24845 6392 -20455 6420
rect -24845 6320 -20575 6392
rect -24845 2320 -24745 6320
rect -20745 2320 -20575 6320
rect -24845 2248 -20575 2320
rect -20475 2248 -20455 6392
rect -24845 2220 -20455 2248
rect -20315 6392 -15925 6420
rect -20315 6320 -16045 6392
rect -20315 2320 -20215 6320
rect -16215 2320 -16045 6320
rect -20315 2248 -16045 2320
rect -15945 2248 -15925 6392
rect -20315 2220 -15925 2248
rect -15785 6392 -11395 6420
rect -15785 6320 -11515 6392
rect -15785 2320 -15685 6320
rect -11685 2320 -11515 6320
rect -15785 2248 -11515 2320
rect -11415 2248 -11395 6392
rect -15785 2220 -11395 2248
rect -11255 6392 -6865 6420
rect -11255 6320 -6985 6392
rect -11255 2320 -11155 6320
rect -7155 2320 -6985 6320
rect -11255 2248 -6985 2320
rect -6885 2248 -6865 6392
rect -11255 2220 -6865 2248
rect -6725 6392 -2335 6420
rect -6725 6320 -2455 6392
rect -6725 2320 -6625 6320
rect -2625 2320 -2455 6320
rect -6725 2248 -2455 2320
rect -2355 2248 -2335 6392
rect -6725 2220 -2335 2248
rect -2195 6392 2195 6420
rect -2195 6320 2075 6392
rect -2195 2320 -2095 6320
rect 1905 2320 2075 6320
rect -2195 2248 2075 2320
rect 2175 2248 2195 6392
rect -2195 2220 2195 2248
rect 2335 6392 6725 6420
rect 2335 6320 6605 6392
rect 2335 2320 2435 6320
rect 6435 2320 6605 6320
rect 2335 2248 6605 2320
rect 6705 2248 6725 6392
rect 2335 2220 6725 2248
rect 6865 6392 11255 6420
rect 6865 6320 11135 6392
rect 6865 2320 6965 6320
rect 10965 2320 11135 6320
rect 6865 2248 11135 2320
rect 11235 2248 11255 6392
rect 6865 2220 11255 2248
rect 11395 6392 15785 6420
rect 11395 6320 15665 6392
rect 11395 2320 11495 6320
rect 15495 2320 15665 6320
rect 11395 2248 15665 2320
rect 15765 2248 15785 6392
rect 11395 2220 15785 2248
rect 15925 6392 20315 6420
rect 15925 6320 20195 6392
rect 15925 2320 16025 6320
rect 20025 2320 20195 6320
rect 15925 2248 20195 2320
rect 20295 2248 20315 6392
rect 15925 2220 20315 2248
rect 20455 6392 24845 6420
rect 20455 6320 24725 6392
rect 20455 2320 20555 6320
rect 24555 2320 24725 6320
rect 20455 2248 24725 2320
rect 24825 2248 24845 6392
rect 20455 2220 24845 2248
rect 24985 6392 29375 6420
rect 24985 6320 29255 6392
rect 24985 2320 25085 6320
rect 29085 2320 29255 6320
rect 24985 2248 29255 2320
rect 29355 2248 29375 6392
rect 24985 2220 29375 2248
rect 29515 6392 33905 6420
rect 29515 6320 33785 6392
rect 29515 2320 29615 6320
rect 33615 2320 33785 6320
rect 29515 2248 33785 2320
rect 33885 2248 33905 6392
rect 29515 2220 33905 2248
rect 34045 6392 38435 6420
rect 34045 6320 38315 6392
rect 34045 2320 34145 6320
rect 38145 2320 38315 6320
rect 34045 2248 38315 2320
rect 38415 2248 38435 6392
rect 34045 2220 38435 2248
rect 38575 6392 42965 6420
rect 38575 6320 42845 6392
rect 38575 2320 38675 6320
rect 42675 2320 42845 6320
rect 38575 2248 42845 2320
rect 42945 2248 42965 6392
rect 38575 2220 42965 2248
rect 43105 6392 47495 6420
rect 43105 6320 47375 6392
rect 43105 2320 43205 6320
rect 47205 2320 47375 6320
rect 43105 2248 47375 2320
rect 47475 2248 47495 6392
rect 43105 2220 47495 2248
rect 47635 6392 52025 6420
rect 47635 6320 51905 6392
rect 47635 2320 47735 6320
rect 51735 2320 51905 6320
rect 47635 2248 51905 2320
rect 52005 2248 52025 6392
rect 47635 2220 52025 2248
rect 52165 6392 56555 6420
rect 52165 6320 56435 6392
rect 52165 2320 52265 6320
rect 56265 2320 56435 6320
rect 52165 2248 56435 2320
rect 56535 2248 56555 6392
rect 52165 2220 56555 2248
rect 56695 6392 61085 6420
rect 56695 6320 60965 6392
rect 56695 2320 56795 6320
rect 60795 2320 60965 6320
rect 56695 2248 60965 2320
rect 61065 2248 61085 6392
rect 56695 2220 61085 2248
rect 61225 6392 65615 6420
rect 61225 6320 65495 6392
rect 61225 2320 61325 6320
rect 65325 2320 65495 6320
rect 61225 2248 65495 2320
rect 65595 2248 65615 6392
rect 61225 2220 65615 2248
rect 65755 6392 70145 6420
rect 65755 6320 70025 6392
rect 65755 2320 65855 6320
rect 69855 2320 70025 6320
rect 65755 2248 70025 2320
rect 70125 2248 70145 6392
rect 65755 2220 70145 2248
rect 70285 6392 74675 6420
rect 70285 6320 74555 6392
rect 70285 2320 70385 6320
rect 74385 2320 74555 6320
rect 70285 2248 74555 2320
rect 74655 2248 74675 6392
rect 70285 2220 74675 2248
rect 74815 6392 79205 6420
rect 74815 6320 79085 6392
rect 74815 2320 74915 6320
rect 78915 2320 79085 6320
rect 74815 2248 79085 2320
rect 79185 2248 79205 6392
rect 74815 2220 79205 2248
rect 79345 6392 83735 6420
rect 79345 6320 83615 6392
rect 79345 2320 79445 6320
rect 83445 2320 83615 6320
rect 79345 2248 83615 2320
rect 83715 2248 83735 6392
rect 79345 2220 83735 2248
rect 83875 6392 88265 6420
rect 83875 6320 88145 6392
rect 83875 2320 83975 6320
rect 87975 2320 88145 6320
rect 83875 2248 88145 2320
rect 88245 2248 88265 6392
rect 83875 2220 88265 2248
rect 88405 6392 92795 6420
rect 88405 6320 92675 6392
rect 88405 2320 88505 6320
rect 92505 2320 92675 6320
rect 88405 2248 92675 2320
rect 92775 2248 92795 6392
rect 88405 2220 92795 2248
rect 92935 6392 97325 6420
rect 92935 6320 97205 6392
rect 92935 2320 93035 6320
rect 97035 2320 97205 6320
rect 92935 2248 97205 2320
rect 97305 2248 97325 6392
rect 92935 2220 97325 2248
rect 97465 6392 101855 6420
rect 97465 6320 101735 6392
rect 97465 2320 97565 6320
rect 101565 2320 101735 6320
rect 97465 2248 101735 2320
rect 101835 2248 101855 6392
rect 97465 2220 101855 2248
rect 101995 6392 106385 6420
rect 101995 6320 106265 6392
rect 101995 2320 102095 6320
rect 106095 2320 106265 6320
rect 101995 2248 106265 2320
rect 106365 2248 106385 6392
rect 101995 2220 106385 2248
rect 106525 6392 110915 6420
rect 106525 6320 110795 6392
rect 106525 2320 106625 6320
rect 110625 2320 110795 6320
rect 106525 2248 110795 2320
rect 110895 2248 110915 6392
rect 106525 2220 110915 2248
rect 111055 6392 115445 6420
rect 111055 6320 115325 6392
rect 111055 2320 111155 6320
rect 115155 2320 115325 6320
rect 111055 2248 115325 2320
rect 115425 2248 115445 6392
rect 111055 2220 115445 2248
rect 115585 6392 119975 6420
rect 115585 6320 119855 6392
rect 115585 2320 115685 6320
rect 119685 2320 119855 6320
rect 115585 2248 119855 2320
rect 119955 2248 119975 6392
rect 115585 2220 119975 2248
rect 120115 6392 124505 6420
rect 120115 6320 124385 6392
rect 120115 2320 120215 6320
rect 124215 2320 124385 6320
rect 120115 2248 124385 2320
rect 124485 2248 124505 6392
rect 120115 2220 124505 2248
rect -124505 2072 -120115 2100
rect -124505 2000 -120235 2072
rect -124505 -2000 -124405 2000
rect -120405 -2000 -120235 2000
rect -124505 -2072 -120235 -2000
rect -120135 -2072 -120115 2072
rect -124505 -2100 -120115 -2072
rect -119975 2072 -115585 2100
rect -119975 2000 -115705 2072
rect -119975 -2000 -119875 2000
rect -115875 -2000 -115705 2000
rect -119975 -2072 -115705 -2000
rect -115605 -2072 -115585 2072
rect -119975 -2100 -115585 -2072
rect -115445 2072 -111055 2100
rect -115445 2000 -111175 2072
rect -115445 -2000 -115345 2000
rect -111345 -2000 -111175 2000
rect -115445 -2072 -111175 -2000
rect -111075 -2072 -111055 2072
rect -115445 -2100 -111055 -2072
rect -110915 2072 -106525 2100
rect -110915 2000 -106645 2072
rect -110915 -2000 -110815 2000
rect -106815 -2000 -106645 2000
rect -110915 -2072 -106645 -2000
rect -106545 -2072 -106525 2072
rect -110915 -2100 -106525 -2072
rect -106385 2072 -101995 2100
rect -106385 2000 -102115 2072
rect -106385 -2000 -106285 2000
rect -102285 -2000 -102115 2000
rect -106385 -2072 -102115 -2000
rect -102015 -2072 -101995 2072
rect -106385 -2100 -101995 -2072
rect -101855 2072 -97465 2100
rect -101855 2000 -97585 2072
rect -101855 -2000 -101755 2000
rect -97755 -2000 -97585 2000
rect -101855 -2072 -97585 -2000
rect -97485 -2072 -97465 2072
rect -101855 -2100 -97465 -2072
rect -97325 2072 -92935 2100
rect -97325 2000 -93055 2072
rect -97325 -2000 -97225 2000
rect -93225 -2000 -93055 2000
rect -97325 -2072 -93055 -2000
rect -92955 -2072 -92935 2072
rect -97325 -2100 -92935 -2072
rect -92795 2072 -88405 2100
rect -92795 2000 -88525 2072
rect -92795 -2000 -92695 2000
rect -88695 -2000 -88525 2000
rect -92795 -2072 -88525 -2000
rect -88425 -2072 -88405 2072
rect -92795 -2100 -88405 -2072
rect -88265 2072 -83875 2100
rect -88265 2000 -83995 2072
rect -88265 -2000 -88165 2000
rect -84165 -2000 -83995 2000
rect -88265 -2072 -83995 -2000
rect -83895 -2072 -83875 2072
rect -88265 -2100 -83875 -2072
rect -83735 2072 -79345 2100
rect -83735 2000 -79465 2072
rect -83735 -2000 -83635 2000
rect -79635 -2000 -79465 2000
rect -83735 -2072 -79465 -2000
rect -79365 -2072 -79345 2072
rect -83735 -2100 -79345 -2072
rect -79205 2072 -74815 2100
rect -79205 2000 -74935 2072
rect -79205 -2000 -79105 2000
rect -75105 -2000 -74935 2000
rect -79205 -2072 -74935 -2000
rect -74835 -2072 -74815 2072
rect -79205 -2100 -74815 -2072
rect -74675 2072 -70285 2100
rect -74675 2000 -70405 2072
rect -74675 -2000 -74575 2000
rect -70575 -2000 -70405 2000
rect -74675 -2072 -70405 -2000
rect -70305 -2072 -70285 2072
rect -74675 -2100 -70285 -2072
rect -70145 2072 -65755 2100
rect -70145 2000 -65875 2072
rect -70145 -2000 -70045 2000
rect -66045 -2000 -65875 2000
rect -70145 -2072 -65875 -2000
rect -65775 -2072 -65755 2072
rect -70145 -2100 -65755 -2072
rect -65615 2072 -61225 2100
rect -65615 2000 -61345 2072
rect -65615 -2000 -65515 2000
rect -61515 -2000 -61345 2000
rect -65615 -2072 -61345 -2000
rect -61245 -2072 -61225 2072
rect -65615 -2100 -61225 -2072
rect -61085 2072 -56695 2100
rect -61085 2000 -56815 2072
rect -61085 -2000 -60985 2000
rect -56985 -2000 -56815 2000
rect -61085 -2072 -56815 -2000
rect -56715 -2072 -56695 2072
rect -61085 -2100 -56695 -2072
rect -56555 2072 -52165 2100
rect -56555 2000 -52285 2072
rect -56555 -2000 -56455 2000
rect -52455 -2000 -52285 2000
rect -56555 -2072 -52285 -2000
rect -52185 -2072 -52165 2072
rect -56555 -2100 -52165 -2072
rect -52025 2072 -47635 2100
rect -52025 2000 -47755 2072
rect -52025 -2000 -51925 2000
rect -47925 -2000 -47755 2000
rect -52025 -2072 -47755 -2000
rect -47655 -2072 -47635 2072
rect -52025 -2100 -47635 -2072
rect -47495 2072 -43105 2100
rect -47495 2000 -43225 2072
rect -47495 -2000 -47395 2000
rect -43395 -2000 -43225 2000
rect -47495 -2072 -43225 -2000
rect -43125 -2072 -43105 2072
rect -47495 -2100 -43105 -2072
rect -42965 2072 -38575 2100
rect -42965 2000 -38695 2072
rect -42965 -2000 -42865 2000
rect -38865 -2000 -38695 2000
rect -42965 -2072 -38695 -2000
rect -38595 -2072 -38575 2072
rect -42965 -2100 -38575 -2072
rect -38435 2072 -34045 2100
rect -38435 2000 -34165 2072
rect -38435 -2000 -38335 2000
rect -34335 -2000 -34165 2000
rect -38435 -2072 -34165 -2000
rect -34065 -2072 -34045 2072
rect -38435 -2100 -34045 -2072
rect -33905 2072 -29515 2100
rect -33905 2000 -29635 2072
rect -33905 -2000 -33805 2000
rect -29805 -2000 -29635 2000
rect -33905 -2072 -29635 -2000
rect -29535 -2072 -29515 2072
rect -33905 -2100 -29515 -2072
rect -29375 2072 -24985 2100
rect -29375 2000 -25105 2072
rect -29375 -2000 -29275 2000
rect -25275 -2000 -25105 2000
rect -29375 -2072 -25105 -2000
rect -25005 -2072 -24985 2072
rect -29375 -2100 -24985 -2072
rect -24845 2072 -20455 2100
rect -24845 2000 -20575 2072
rect -24845 -2000 -24745 2000
rect -20745 -2000 -20575 2000
rect -24845 -2072 -20575 -2000
rect -20475 -2072 -20455 2072
rect -24845 -2100 -20455 -2072
rect -20315 2072 -15925 2100
rect -20315 2000 -16045 2072
rect -20315 -2000 -20215 2000
rect -16215 -2000 -16045 2000
rect -20315 -2072 -16045 -2000
rect -15945 -2072 -15925 2072
rect -20315 -2100 -15925 -2072
rect -15785 2072 -11395 2100
rect -15785 2000 -11515 2072
rect -15785 -2000 -15685 2000
rect -11685 -2000 -11515 2000
rect -15785 -2072 -11515 -2000
rect -11415 -2072 -11395 2072
rect -15785 -2100 -11395 -2072
rect -11255 2072 -6865 2100
rect -11255 2000 -6985 2072
rect -11255 -2000 -11155 2000
rect -7155 -2000 -6985 2000
rect -11255 -2072 -6985 -2000
rect -6885 -2072 -6865 2072
rect -11255 -2100 -6865 -2072
rect -6725 2072 -2335 2100
rect -6725 2000 -2455 2072
rect -6725 -2000 -6625 2000
rect -2625 -2000 -2455 2000
rect -6725 -2072 -2455 -2000
rect -2355 -2072 -2335 2072
rect -6725 -2100 -2335 -2072
rect -2195 2072 2195 2100
rect -2195 2000 2075 2072
rect -2195 -2000 -2095 2000
rect 1905 -2000 2075 2000
rect -2195 -2072 2075 -2000
rect 2175 -2072 2195 2072
rect -2195 -2100 2195 -2072
rect 2335 2072 6725 2100
rect 2335 2000 6605 2072
rect 2335 -2000 2435 2000
rect 6435 -2000 6605 2000
rect 2335 -2072 6605 -2000
rect 6705 -2072 6725 2072
rect 2335 -2100 6725 -2072
rect 6865 2072 11255 2100
rect 6865 2000 11135 2072
rect 6865 -2000 6965 2000
rect 10965 -2000 11135 2000
rect 6865 -2072 11135 -2000
rect 11235 -2072 11255 2072
rect 6865 -2100 11255 -2072
rect 11395 2072 15785 2100
rect 11395 2000 15665 2072
rect 11395 -2000 11495 2000
rect 15495 -2000 15665 2000
rect 11395 -2072 15665 -2000
rect 15765 -2072 15785 2072
rect 11395 -2100 15785 -2072
rect 15925 2072 20315 2100
rect 15925 2000 20195 2072
rect 15925 -2000 16025 2000
rect 20025 -2000 20195 2000
rect 15925 -2072 20195 -2000
rect 20295 -2072 20315 2072
rect 15925 -2100 20315 -2072
rect 20455 2072 24845 2100
rect 20455 2000 24725 2072
rect 20455 -2000 20555 2000
rect 24555 -2000 24725 2000
rect 20455 -2072 24725 -2000
rect 24825 -2072 24845 2072
rect 20455 -2100 24845 -2072
rect 24985 2072 29375 2100
rect 24985 2000 29255 2072
rect 24985 -2000 25085 2000
rect 29085 -2000 29255 2000
rect 24985 -2072 29255 -2000
rect 29355 -2072 29375 2072
rect 24985 -2100 29375 -2072
rect 29515 2072 33905 2100
rect 29515 2000 33785 2072
rect 29515 -2000 29615 2000
rect 33615 -2000 33785 2000
rect 29515 -2072 33785 -2000
rect 33885 -2072 33905 2072
rect 29515 -2100 33905 -2072
rect 34045 2072 38435 2100
rect 34045 2000 38315 2072
rect 34045 -2000 34145 2000
rect 38145 -2000 38315 2000
rect 34045 -2072 38315 -2000
rect 38415 -2072 38435 2072
rect 34045 -2100 38435 -2072
rect 38575 2072 42965 2100
rect 38575 2000 42845 2072
rect 38575 -2000 38675 2000
rect 42675 -2000 42845 2000
rect 38575 -2072 42845 -2000
rect 42945 -2072 42965 2072
rect 38575 -2100 42965 -2072
rect 43105 2072 47495 2100
rect 43105 2000 47375 2072
rect 43105 -2000 43205 2000
rect 47205 -2000 47375 2000
rect 43105 -2072 47375 -2000
rect 47475 -2072 47495 2072
rect 43105 -2100 47495 -2072
rect 47635 2072 52025 2100
rect 47635 2000 51905 2072
rect 47635 -2000 47735 2000
rect 51735 -2000 51905 2000
rect 47635 -2072 51905 -2000
rect 52005 -2072 52025 2072
rect 47635 -2100 52025 -2072
rect 52165 2072 56555 2100
rect 52165 2000 56435 2072
rect 52165 -2000 52265 2000
rect 56265 -2000 56435 2000
rect 52165 -2072 56435 -2000
rect 56535 -2072 56555 2072
rect 52165 -2100 56555 -2072
rect 56695 2072 61085 2100
rect 56695 2000 60965 2072
rect 56695 -2000 56795 2000
rect 60795 -2000 60965 2000
rect 56695 -2072 60965 -2000
rect 61065 -2072 61085 2072
rect 56695 -2100 61085 -2072
rect 61225 2072 65615 2100
rect 61225 2000 65495 2072
rect 61225 -2000 61325 2000
rect 65325 -2000 65495 2000
rect 61225 -2072 65495 -2000
rect 65595 -2072 65615 2072
rect 61225 -2100 65615 -2072
rect 65755 2072 70145 2100
rect 65755 2000 70025 2072
rect 65755 -2000 65855 2000
rect 69855 -2000 70025 2000
rect 65755 -2072 70025 -2000
rect 70125 -2072 70145 2072
rect 65755 -2100 70145 -2072
rect 70285 2072 74675 2100
rect 70285 2000 74555 2072
rect 70285 -2000 70385 2000
rect 74385 -2000 74555 2000
rect 70285 -2072 74555 -2000
rect 74655 -2072 74675 2072
rect 70285 -2100 74675 -2072
rect 74815 2072 79205 2100
rect 74815 2000 79085 2072
rect 74815 -2000 74915 2000
rect 78915 -2000 79085 2000
rect 74815 -2072 79085 -2000
rect 79185 -2072 79205 2072
rect 74815 -2100 79205 -2072
rect 79345 2072 83735 2100
rect 79345 2000 83615 2072
rect 79345 -2000 79445 2000
rect 83445 -2000 83615 2000
rect 79345 -2072 83615 -2000
rect 83715 -2072 83735 2072
rect 79345 -2100 83735 -2072
rect 83875 2072 88265 2100
rect 83875 2000 88145 2072
rect 83875 -2000 83975 2000
rect 87975 -2000 88145 2000
rect 83875 -2072 88145 -2000
rect 88245 -2072 88265 2072
rect 83875 -2100 88265 -2072
rect 88405 2072 92795 2100
rect 88405 2000 92675 2072
rect 88405 -2000 88505 2000
rect 92505 -2000 92675 2000
rect 88405 -2072 92675 -2000
rect 92775 -2072 92795 2072
rect 88405 -2100 92795 -2072
rect 92935 2072 97325 2100
rect 92935 2000 97205 2072
rect 92935 -2000 93035 2000
rect 97035 -2000 97205 2000
rect 92935 -2072 97205 -2000
rect 97305 -2072 97325 2072
rect 92935 -2100 97325 -2072
rect 97465 2072 101855 2100
rect 97465 2000 101735 2072
rect 97465 -2000 97565 2000
rect 101565 -2000 101735 2000
rect 97465 -2072 101735 -2000
rect 101835 -2072 101855 2072
rect 97465 -2100 101855 -2072
rect 101995 2072 106385 2100
rect 101995 2000 106265 2072
rect 101995 -2000 102095 2000
rect 106095 -2000 106265 2000
rect 101995 -2072 106265 -2000
rect 106365 -2072 106385 2072
rect 101995 -2100 106385 -2072
rect 106525 2072 110915 2100
rect 106525 2000 110795 2072
rect 106525 -2000 106625 2000
rect 110625 -2000 110795 2000
rect 106525 -2072 110795 -2000
rect 110895 -2072 110915 2072
rect 106525 -2100 110915 -2072
rect 111055 2072 115445 2100
rect 111055 2000 115325 2072
rect 111055 -2000 111155 2000
rect 115155 -2000 115325 2000
rect 111055 -2072 115325 -2000
rect 115425 -2072 115445 2072
rect 111055 -2100 115445 -2072
rect 115585 2072 119975 2100
rect 115585 2000 119855 2072
rect 115585 -2000 115685 2000
rect 119685 -2000 119855 2000
rect 115585 -2072 119855 -2000
rect 119955 -2072 119975 2072
rect 115585 -2100 119975 -2072
rect 120115 2072 124505 2100
rect 120115 2000 124385 2072
rect 120115 -2000 120215 2000
rect 124215 -2000 124385 2000
rect 120115 -2072 124385 -2000
rect 124485 -2072 124505 2072
rect 120115 -2100 124505 -2072
rect -124505 -2248 -120115 -2220
rect -124505 -2320 -120235 -2248
rect -124505 -6320 -124405 -2320
rect -120405 -6320 -120235 -2320
rect -124505 -6392 -120235 -6320
rect -120135 -6392 -120115 -2248
rect -124505 -6420 -120115 -6392
rect -119975 -2248 -115585 -2220
rect -119975 -2320 -115705 -2248
rect -119975 -6320 -119875 -2320
rect -115875 -6320 -115705 -2320
rect -119975 -6392 -115705 -6320
rect -115605 -6392 -115585 -2248
rect -119975 -6420 -115585 -6392
rect -115445 -2248 -111055 -2220
rect -115445 -2320 -111175 -2248
rect -115445 -6320 -115345 -2320
rect -111345 -6320 -111175 -2320
rect -115445 -6392 -111175 -6320
rect -111075 -6392 -111055 -2248
rect -115445 -6420 -111055 -6392
rect -110915 -2248 -106525 -2220
rect -110915 -2320 -106645 -2248
rect -110915 -6320 -110815 -2320
rect -106815 -6320 -106645 -2320
rect -110915 -6392 -106645 -6320
rect -106545 -6392 -106525 -2248
rect -110915 -6420 -106525 -6392
rect -106385 -2248 -101995 -2220
rect -106385 -2320 -102115 -2248
rect -106385 -6320 -106285 -2320
rect -102285 -6320 -102115 -2320
rect -106385 -6392 -102115 -6320
rect -102015 -6392 -101995 -2248
rect -106385 -6420 -101995 -6392
rect -101855 -2248 -97465 -2220
rect -101855 -2320 -97585 -2248
rect -101855 -6320 -101755 -2320
rect -97755 -6320 -97585 -2320
rect -101855 -6392 -97585 -6320
rect -97485 -6392 -97465 -2248
rect -101855 -6420 -97465 -6392
rect -97325 -2248 -92935 -2220
rect -97325 -2320 -93055 -2248
rect -97325 -6320 -97225 -2320
rect -93225 -6320 -93055 -2320
rect -97325 -6392 -93055 -6320
rect -92955 -6392 -92935 -2248
rect -97325 -6420 -92935 -6392
rect -92795 -2248 -88405 -2220
rect -92795 -2320 -88525 -2248
rect -92795 -6320 -92695 -2320
rect -88695 -6320 -88525 -2320
rect -92795 -6392 -88525 -6320
rect -88425 -6392 -88405 -2248
rect -92795 -6420 -88405 -6392
rect -88265 -2248 -83875 -2220
rect -88265 -2320 -83995 -2248
rect -88265 -6320 -88165 -2320
rect -84165 -6320 -83995 -2320
rect -88265 -6392 -83995 -6320
rect -83895 -6392 -83875 -2248
rect -88265 -6420 -83875 -6392
rect -83735 -2248 -79345 -2220
rect -83735 -2320 -79465 -2248
rect -83735 -6320 -83635 -2320
rect -79635 -6320 -79465 -2320
rect -83735 -6392 -79465 -6320
rect -79365 -6392 -79345 -2248
rect -83735 -6420 -79345 -6392
rect -79205 -2248 -74815 -2220
rect -79205 -2320 -74935 -2248
rect -79205 -6320 -79105 -2320
rect -75105 -6320 -74935 -2320
rect -79205 -6392 -74935 -6320
rect -74835 -6392 -74815 -2248
rect -79205 -6420 -74815 -6392
rect -74675 -2248 -70285 -2220
rect -74675 -2320 -70405 -2248
rect -74675 -6320 -74575 -2320
rect -70575 -6320 -70405 -2320
rect -74675 -6392 -70405 -6320
rect -70305 -6392 -70285 -2248
rect -74675 -6420 -70285 -6392
rect -70145 -2248 -65755 -2220
rect -70145 -2320 -65875 -2248
rect -70145 -6320 -70045 -2320
rect -66045 -6320 -65875 -2320
rect -70145 -6392 -65875 -6320
rect -65775 -6392 -65755 -2248
rect -70145 -6420 -65755 -6392
rect -65615 -2248 -61225 -2220
rect -65615 -2320 -61345 -2248
rect -65615 -6320 -65515 -2320
rect -61515 -6320 -61345 -2320
rect -65615 -6392 -61345 -6320
rect -61245 -6392 -61225 -2248
rect -65615 -6420 -61225 -6392
rect -61085 -2248 -56695 -2220
rect -61085 -2320 -56815 -2248
rect -61085 -6320 -60985 -2320
rect -56985 -6320 -56815 -2320
rect -61085 -6392 -56815 -6320
rect -56715 -6392 -56695 -2248
rect -61085 -6420 -56695 -6392
rect -56555 -2248 -52165 -2220
rect -56555 -2320 -52285 -2248
rect -56555 -6320 -56455 -2320
rect -52455 -6320 -52285 -2320
rect -56555 -6392 -52285 -6320
rect -52185 -6392 -52165 -2248
rect -56555 -6420 -52165 -6392
rect -52025 -2248 -47635 -2220
rect -52025 -2320 -47755 -2248
rect -52025 -6320 -51925 -2320
rect -47925 -6320 -47755 -2320
rect -52025 -6392 -47755 -6320
rect -47655 -6392 -47635 -2248
rect -52025 -6420 -47635 -6392
rect -47495 -2248 -43105 -2220
rect -47495 -2320 -43225 -2248
rect -47495 -6320 -47395 -2320
rect -43395 -6320 -43225 -2320
rect -47495 -6392 -43225 -6320
rect -43125 -6392 -43105 -2248
rect -47495 -6420 -43105 -6392
rect -42965 -2248 -38575 -2220
rect -42965 -2320 -38695 -2248
rect -42965 -6320 -42865 -2320
rect -38865 -6320 -38695 -2320
rect -42965 -6392 -38695 -6320
rect -38595 -6392 -38575 -2248
rect -42965 -6420 -38575 -6392
rect -38435 -2248 -34045 -2220
rect -38435 -2320 -34165 -2248
rect -38435 -6320 -38335 -2320
rect -34335 -6320 -34165 -2320
rect -38435 -6392 -34165 -6320
rect -34065 -6392 -34045 -2248
rect -38435 -6420 -34045 -6392
rect -33905 -2248 -29515 -2220
rect -33905 -2320 -29635 -2248
rect -33905 -6320 -33805 -2320
rect -29805 -6320 -29635 -2320
rect -33905 -6392 -29635 -6320
rect -29535 -6392 -29515 -2248
rect -33905 -6420 -29515 -6392
rect -29375 -2248 -24985 -2220
rect -29375 -2320 -25105 -2248
rect -29375 -6320 -29275 -2320
rect -25275 -6320 -25105 -2320
rect -29375 -6392 -25105 -6320
rect -25005 -6392 -24985 -2248
rect -29375 -6420 -24985 -6392
rect -24845 -2248 -20455 -2220
rect -24845 -2320 -20575 -2248
rect -24845 -6320 -24745 -2320
rect -20745 -6320 -20575 -2320
rect -24845 -6392 -20575 -6320
rect -20475 -6392 -20455 -2248
rect -24845 -6420 -20455 -6392
rect -20315 -2248 -15925 -2220
rect -20315 -2320 -16045 -2248
rect -20315 -6320 -20215 -2320
rect -16215 -6320 -16045 -2320
rect -20315 -6392 -16045 -6320
rect -15945 -6392 -15925 -2248
rect -20315 -6420 -15925 -6392
rect -15785 -2248 -11395 -2220
rect -15785 -2320 -11515 -2248
rect -15785 -6320 -15685 -2320
rect -11685 -6320 -11515 -2320
rect -15785 -6392 -11515 -6320
rect -11415 -6392 -11395 -2248
rect -15785 -6420 -11395 -6392
rect -11255 -2248 -6865 -2220
rect -11255 -2320 -6985 -2248
rect -11255 -6320 -11155 -2320
rect -7155 -6320 -6985 -2320
rect -11255 -6392 -6985 -6320
rect -6885 -6392 -6865 -2248
rect -11255 -6420 -6865 -6392
rect -6725 -2248 -2335 -2220
rect -6725 -2320 -2455 -2248
rect -6725 -6320 -6625 -2320
rect -2625 -6320 -2455 -2320
rect -6725 -6392 -2455 -6320
rect -2355 -6392 -2335 -2248
rect -6725 -6420 -2335 -6392
rect -2195 -2248 2195 -2220
rect -2195 -2320 2075 -2248
rect -2195 -6320 -2095 -2320
rect 1905 -6320 2075 -2320
rect -2195 -6392 2075 -6320
rect 2175 -6392 2195 -2248
rect -2195 -6420 2195 -6392
rect 2335 -2248 6725 -2220
rect 2335 -2320 6605 -2248
rect 2335 -6320 2435 -2320
rect 6435 -6320 6605 -2320
rect 2335 -6392 6605 -6320
rect 6705 -6392 6725 -2248
rect 2335 -6420 6725 -6392
rect 6865 -2248 11255 -2220
rect 6865 -2320 11135 -2248
rect 6865 -6320 6965 -2320
rect 10965 -6320 11135 -2320
rect 6865 -6392 11135 -6320
rect 11235 -6392 11255 -2248
rect 6865 -6420 11255 -6392
rect 11395 -2248 15785 -2220
rect 11395 -2320 15665 -2248
rect 11395 -6320 11495 -2320
rect 15495 -6320 15665 -2320
rect 11395 -6392 15665 -6320
rect 15765 -6392 15785 -2248
rect 11395 -6420 15785 -6392
rect 15925 -2248 20315 -2220
rect 15925 -2320 20195 -2248
rect 15925 -6320 16025 -2320
rect 20025 -6320 20195 -2320
rect 15925 -6392 20195 -6320
rect 20295 -6392 20315 -2248
rect 15925 -6420 20315 -6392
rect 20455 -2248 24845 -2220
rect 20455 -2320 24725 -2248
rect 20455 -6320 20555 -2320
rect 24555 -6320 24725 -2320
rect 20455 -6392 24725 -6320
rect 24825 -6392 24845 -2248
rect 20455 -6420 24845 -6392
rect 24985 -2248 29375 -2220
rect 24985 -2320 29255 -2248
rect 24985 -6320 25085 -2320
rect 29085 -6320 29255 -2320
rect 24985 -6392 29255 -6320
rect 29355 -6392 29375 -2248
rect 24985 -6420 29375 -6392
rect 29515 -2248 33905 -2220
rect 29515 -2320 33785 -2248
rect 29515 -6320 29615 -2320
rect 33615 -6320 33785 -2320
rect 29515 -6392 33785 -6320
rect 33885 -6392 33905 -2248
rect 29515 -6420 33905 -6392
rect 34045 -2248 38435 -2220
rect 34045 -2320 38315 -2248
rect 34045 -6320 34145 -2320
rect 38145 -6320 38315 -2320
rect 34045 -6392 38315 -6320
rect 38415 -6392 38435 -2248
rect 34045 -6420 38435 -6392
rect 38575 -2248 42965 -2220
rect 38575 -2320 42845 -2248
rect 38575 -6320 38675 -2320
rect 42675 -6320 42845 -2320
rect 38575 -6392 42845 -6320
rect 42945 -6392 42965 -2248
rect 38575 -6420 42965 -6392
rect 43105 -2248 47495 -2220
rect 43105 -2320 47375 -2248
rect 43105 -6320 43205 -2320
rect 47205 -6320 47375 -2320
rect 43105 -6392 47375 -6320
rect 47475 -6392 47495 -2248
rect 43105 -6420 47495 -6392
rect 47635 -2248 52025 -2220
rect 47635 -2320 51905 -2248
rect 47635 -6320 47735 -2320
rect 51735 -6320 51905 -2320
rect 47635 -6392 51905 -6320
rect 52005 -6392 52025 -2248
rect 47635 -6420 52025 -6392
rect 52165 -2248 56555 -2220
rect 52165 -2320 56435 -2248
rect 52165 -6320 52265 -2320
rect 56265 -6320 56435 -2320
rect 52165 -6392 56435 -6320
rect 56535 -6392 56555 -2248
rect 52165 -6420 56555 -6392
rect 56695 -2248 61085 -2220
rect 56695 -2320 60965 -2248
rect 56695 -6320 56795 -2320
rect 60795 -6320 60965 -2320
rect 56695 -6392 60965 -6320
rect 61065 -6392 61085 -2248
rect 56695 -6420 61085 -6392
rect 61225 -2248 65615 -2220
rect 61225 -2320 65495 -2248
rect 61225 -6320 61325 -2320
rect 65325 -6320 65495 -2320
rect 61225 -6392 65495 -6320
rect 65595 -6392 65615 -2248
rect 61225 -6420 65615 -6392
rect 65755 -2248 70145 -2220
rect 65755 -2320 70025 -2248
rect 65755 -6320 65855 -2320
rect 69855 -6320 70025 -2320
rect 65755 -6392 70025 -6320
rect 70125 -6392 70145 -2248
rect 65755 -6420 70145 -6392
rect 70285 -2248 74675 -2220
rect 70285 -2320 74555 -2248
rect 70285 -6320 70385 -2320
rect 74385 -6320 74555 -2320
rect 70285 -6392 74555 -6320
rect 74655 -6392 74675 -2248
rect 70285 -6420 74675 -6392
rect 74815 -2248 79205 -2220
rect 74815 -2320 79085 -2248
rect 74815 -6320 74915 -2320
rect 78915 -6320 79085 -2320
rect 74815 -6392 79085 -6320
rect 79185 -6392 79205 -2248
rect 74815 -6420 79205 -6392
rect 79345 -2248 83735 -2220
rect 79345 -2320 83615 -2248
rect 79345 -6320 79445 -2320
rect 83445 -6320 83615 -2320
rect 79345 -6392 83615 -6320
rect 83715 -6392 83735 -2248
rect 79345 -6420 83735 -6392
rect 83875 -2248 88265 -2220
rect 83875 -2320 88145 -2248
rect 83875 -6320 83975 -2320
rect 87975 -6320 88145 -2320
rect 83875 -6392 88145 -6320
rect 88245 -6392 88265 -2248
rect 83875 -6420 88265 -6392
rect 88405 -2248 92795 -2220
rect 88405 -2320 92675 -2248
rect 88405 -6320 88505 -2320
rect 92505 -6320 92675 -2320
rect 88405 -6392 92675 -6320
rect 92775 -6392 92795 -2248
rect 88405 -6420 92795 -6392
rect 92935 -2248 97325 -2220
rect 92935 -2320 97205 -2248
rect 92935 -6320 93035 -2320
rect 97035 -6320 97205 -2320
rect 92935 -6392 97205 -6320
rect 97305 -6392 97325 -2248
rect 92935 -6420 97325 -6392
rect 97465 -2248 101855 -2220
rect 97465 -2320 101735 -2248
rect 97465 -6320 97565 -2320
rect 101565 -6320 101735 -2320
rect 97465 -6392 101735 -6320
rect 101835 -6392 101855 -2248
rect 97465 -6420 101855 -6392
rect 101995 -2248 106385 -2220
rect 101995 -2320 106265 -2248
rect 101995 -6320 102095 -2320
rect 106095 -6320 106265 -2320
rect 101995 -6392 106265 -6320
rect 106365 -6392 106385 -2248
rect 101995 -6420 106385 -6392
rect 106525 -2248 110915 -2220
rect 106525 -2320 110795 -2248
rect 106525 -6320 106625 -2320
rect 110625 -6320 110795 -2320
rect 106525 -6392 110795 -6320
rect 110895 -6392 110915 -2248
rect 106525 -6420 110915 -6392
rect 111055 -2248 115445 -2220
rect 111055 -2320 115325 -2248
rect 111055 -6320 111155 -2320
rect 115155 -6320 115325 -2320
rect 111055 -6392 115325 -6320
rect 115425 -6392 115445 -2248
rect 111055 -6420 115445 -6392
rect 115585 -2248 119975 -2220
rect 115585 -2320 119855 -2248
rect 115585 -6320 115685 -2320
rect 119685 -6320 119855 -2320
rect 115585 -6392 119855 -6320
rect 119955 -6392 119975 -2248
rect 115585 -6420 119975 -6392
rect 120115 -2248 124505 -2220
rect 120115 -2320 124385 -2248
rect 120115 -6320 120215 -2320
rect 124215 -6320 124385 -2320
rect 120115 -6392 124385 -6320
rect 124485 -6392 124505 -2248
rect 120115 -6420 124505 -6392
<< viatp >>
rect -120235 2248 -120135 6392
rect -115705 2248 -115605 6392
rect -111175 2248 -111075 6392
rect -106645 2248 -106545 6392
rect -102115 2248 -102015 6392
rect -97585 2248 -97485 6392
rect -93055 2248 -92955 6392
rect -88525 2248 -88425 6392
rect -83995 2248 -83895 6392
rect -79465 2248 -79365 6392
rect -74935 2248 -74835 6392
rect -70405 2248 -70305 6392
rect -65875 2248 -65775 6392
rect -61345 2248 -61245 6392
rect -56815 2248 -56715 6392
rect -52285 2248 -52185 6392
rect -47755 2248 -47655 6392
rect -43225 2248 -43125 6392
rect -38695 2248 -38595 6392
rect -34165 2248 -34065 6392
rect -29635 2248 -29535 6392
rect -25105 2248 -25005 6392
rect -20575 2248 -20475 6392
rect -16045 2248 -15945 6392
rect -11515 2248 -11415 6392
rect -6985 2248 -6885 6392
rect -2455 2248 -2355 6392
rect 2075 2248 2175 6392
rect 6605 2248 6705 6392
rect 11135 2248 11235 6392
rect 15665 2248 15765 6392
rect 20195 2248 20295 6392
rect 24725 2248 24825 6392
rect 29255 2248 29355 6392
rect 33785 2248 33885 6392
rect 38315 2248 38415 6392
rect 42845 2248 42945 6392
rect 47375 2248 47475 6392
rect 51905 2248 52005 6392
rect 56435 2248 56535 6392
rect 60965 2248 61065 6392
rect 65495 2248 65595 6392
rect 70025 2248 70125 6392
rect 74555 2248 74655 6392
rect 79085 2248 79185 6392
rect 83615 2248 83715 6392
rect 88145 2248 88245 6392
rect 92675 2248 92775 6392
rect 97205 2248 97305 6392
rect 101735 2248 101835 6392
rect 106265 2248 106365 6392
rect 110795 2248 110895 6392
rect 115325 2248 115425 6392
rect 119855 2248 119955 6392
rect 124385 2248 124485 6392
rect -120235 -2072 -120135 2072
rect -115705 -2072 -115605 2072
rect -111175 -2072 -111075 2072
rect -106645 -2072 -106545 2072
rect -102115 -2072 -102015 2072
rect -97585 -2072 -97485 2072
rect -93055 -2072 -92955 2072
rect -88525 -2072 -88425 2072
rect -83995 -2072 -83895 2072
rect -79465 -2072 -79365 2072
rect -74935 -2072 -74835 2072
rect -70405 -2072 -70305 2072
rect -65875 -2072 -65775 2072
rect -61345 -2072 -61245 2072
rect -56815 -2072 -56715 2072
rect -52285 -2072 -52185 2072
rect -47755 -2072 -47655 2072
rect -43225 -2072 -43125 2072
rect -38695 -2072 -38595 2072
rect -34165 -2072 -34065 2072
rect -29635 -2072 -29535 2072
rect -25105 -2072 -25005 2072
rect -20575 -2072 -20475 2072
rect -16045 -2072 -15945 2072
rect -11515 -2072 -11415 2072
rect -6985 -2072 -6885 2072
rect -2455 -2072 -2355 2072
rect 2075 -2072 2175 2072
rect 6605 -2072 6705 2072
rect 11135 -2072 11235 2072
rect 15665 -2072 15765 2072
rect 20195 -2072 20295 2072
rect 24725 -2072 24825 2072
rect 29255 -2072 29355 2072
rect 33785 -2072 33885 2072
rect 38315 -2072 38415 2072
rect 42845 -2072 42945 2072
rect 47375 -2072 47475 2072
rect 51905 -2072 52005 2072
rect 56435 -2072 56535 2072
rect 60965 -2072 61065 2072
rect 65495 -2072 65595 2072
rect 70025 -2072 70125 2072
rect 74555 -2072 74655 2072
rect 79085 -2072 79185 2072
rect 83615 -2072 83715 2072
rect 88145 -2072 88245 2072
rect 92675 -2072 92775 2072
rect 97205 -2072 97305 2072
rect 101735 -2072 101835 2072
rect 106265 -2072 106365 2072
rect 110795 -2072 110895 2072
rect 115325 -2072 115425 2072
rect 119855 -2072 119955 2072
rect 124385 -2072 124485 2072
rect -120235 -6392 -120135 -2248
rect -115705 -6392 -115605 -2248
rect -111175 -6392 -111075 -2248
rect -106645 -6392 -106545 -2248
rect -102115 -6392 -102015 -2248
rect -97585 -6392 -97485 -2248
rect -93055 -6392 -92955 -2248
rect -88525 -6392 -88425 -2248
rect -83995 -6392 -83895 -2248
rect -79465 -6392 -79365 -2248
rect -74935 -6392 -74835 -2248
rect -70405 -6392 -70305 -2248
rect -65875 -6392 -65775 -2248
rect -61345 -6392 -61245 -2248
rect -56815 -6392 -56715 -2248
rect -52285 -6392 -52185 -2248
rect -47755 -6392 -47655 -2248
rect -43225 -6392 -43125 -2248
rect -38695 -6392 -38595 -2248
rect -34165 -6392 -34065 -2248
rect -29635 -6392 -29535 -2248
rect -25105 -6392 -25005 -2248
rect -20575 -6392 -20475 -2248
rect -16045 -6392 -15945 -2248
rect -11515 -6392 -11415 -2248
rect -6985 -6392 -6885 -2248
rect -2455 -6392 -2355 -2248
rect 2075 -6392 2175 -2248
rect 6605 -6392 6705 -2248
rect 11135 -6392 11235 -2248
rect 15665 -6392 15765 -2248
rect 20195 -6392 20295 -2248
rect 24725 -6392 24825 -2248
rect 29255 -6392 29355 -2248
rect 33785 -6392 33885 -2248
rect 38315 -6392 38415 -2248
rect 42845 -6392 42945 -2248
rect 47375 -6392 47475 -2248
rect 51905 -6392 52005 -2248
rect 56435 -6392 56535 -2248
rect 60965 -6392 61065 -2248
rect 65495 -6392 65595 -2248
rect 70025 -6392 70125 -2248
rect 74555 -6392 74655 -2248
rect 79085 -6392 79185 -2248
rect 83615 -6392 83715 -2248
rect 88145 -6392 88245 -2248
rect 92675 -6392 92775 -2248
rect 97205 -6392 97305 -2248
rect 101735 -6392 101835 -2248
rect 106265 -6392 106365 -2248
rect 110795 -6392 110895 -2248
rect 115325 -6392 115425 -2248
rect 119855 -6392 119955 -2248
rect 124385 -6392 124485 -2248
<< metaltp >>
rect -122475 6290 -122335 6480
rect -120255 6392 -120115 6480
rect -122475 1970 -122335 2350
rect -120255 2248 -120235 6392
rect -120135 2248 -120115 6392
rect -117945 6290 -117805 6480
rect -115725 6392 -115585 6480
rect -120255 2072 -120115 2248
rect -122475 -2350 -122335 -1970
rect -120255 -2072 -120235 2072
rect -120135 -2072 -120115 2072
rect -117945 1970 -117805 2350
rect -115725 2248 -115705 6392
rect -115605 2248 -115585 6392
rect -113415 6290 -113275 6480
rect -111195 6392 -111055 6480
rect -115725 2072 -115585 2248
rect -120255 -2248 -120115 -2072
rect -122475 -6480 -122335 -6290
rect -120255 -6392 -120235 -2248
rect -120135 -6392 -120115 -2248
rect -117945 -2350 -117805 -1970
rect -115725 -2072 -115705 2072
rect -115605 -2072 -115585 2072
rect -113415 1970 -113275 2350
rect -111195 2248 -111175 6392
rect -111075 2248 -111055 6392
rect -108885 6290 -108745 6480
rect -106665 6392 -106525 6480
rect -111195 2072 -111055 2248
rect -115725 -2248 -115585 -2072
rect -120255 -6480 -120115 -6392
rect -117945 -6480 -117805 -6290
rect -115725 -6392 -115705 -2248
rect -115605 -6392 -115585 -2248
rect -113415 -2350 -113275 -1970
rect -111195 -2072 -111175 2072
rect -111075 -2072 -111055 2072
rect -108885 1970 -108745 2350
rect -106665 2248 -106645 6392
rect -106545 2248 -106525 6392
rect -104355 6290 -104215 6480
rect -102135 6392 -101995 6480
rect -106665 2072 -106525 2248
rect -111195 -2248 -111055 -2072
rect -115725 -6480 -115585 -6392
rect -113415 -6480 -113275 -6290
rect -111195 -6392 -111175 -2248
rect -111075 -6392 -111055 -2248
rect -108885 -2350 -108745 -1970
rect -106665 -2072 -106645 2072
rect -106545 -2072 -106525 2072
rect -104355 1970 -104215 2350
rect -102135 2248 -102115 6392
rect -102015 2248 -101995 6392
rect -99825 6290 -99685 6480
rect -97605 6392 -97465 6480
rect -102135 2072 -101995 2248
rect -106665 -2248 -106525 -2072
rect -111195 -6480 -111055 -6392
rect -108885 -6480 -108745 -6290
rect -106665 -6392 -106645 -2248
rect -106545 -6392 -106525 -2248
rect -104355 -2350 -104215 -1970
rect -102135 -2072 -102115 2072
rect -102015 -2072 -101995 2072
rect -99825 1970 -99685 2350
rect -97605 2248 -97585 6392
rect -97485 2248 -97465 6392
rect -95295 6290 -95155 6480
rect -93075 6392 -92935 6480
rect -97605 2072 -97465 2248
rect -102135 -2248 -101995 -2072
rect -106665 -6480 -106525 -6392
rect -104355 -6480 -104215 -6290
rect -102135 -6392 -102115 -2248
rect -102015 -6392 -101995 -2248
rect -99825 -2350 -99685 -1970
rect -97605 -2072 -97585 2072
rect -97485 -2072 -97465 2072
rect -95295 1970 -95155 2350
rect -93075 2248 -93055 6392
rect -92955 2248 -92935 6392
rect -90765 6290 -90625 6480
rect -88545 6392 -88405 6480
rect -93075 2072 -92935 2248
rect -97605 -2248 -97465 -2072
rect -102135 -6480 -101995 -6392
rect -99825 -6480 -99685 -6290
rect -97605 -6392 -97585 -2248
rect -97485 -6392 -97465 -2248
rect -95295 -2350 -95155 -1970
rect -93075 -2072 -93055 2072
rect -92955 -2072 -92935 2072
rect -90765 1970 -90625 2350
rect -88545 2248 -88525 6392
rect -88425 2248 -88405 6392
rect -86235 6290 -86095 6480
rect -84015 6392 -83875 6480
rect -88545 2072 -88405 2248
rect -93075 -2248 -92935 -2072
rect -97605 -6480 -97465 -6392
rect -95295 -6480 -95155 -6290
rect -93075 -6392 -93055 -2248
rect -92955 -6392 -92935 -2248
rect -90765 -2350 -90625 -1970
rect -88545 -2072 -88525 2072
rect -88425 -2072 -88405 2072
rect -86235 1970 -86095 2350
rect -84015 2248 -83995 6392
rect -83895 2248 -83875 6392
rect -81705 6290 -81565 6480
rect -79485 6392 -79345 6480
rect -84015 2072 -83875 2248
rect -88545 -2248 -88405 -2072
rect -93075 -6480 -92935 -6392
rect -90765 -6480 -90625 -6290
rect -88545 -6392 -88525 -2248
rect -88425 -6392 -88405 -2248
rect -86235 -2350 -86095 -1970
rect -84015 -2072 -83995 2072
rect -83895 -2072 -83875 2072
rect -81705 1970 -81565 2350
rect -79485 2248 -79465 6392
rect -79365 2248 -79345 6392
rect -77175 6290 -77035 6480
rect -74955 6392 -74815 6480
rect -79485 2072 -79345 2248
rect -84015 -2248 -83875 -2072
rect -88545 -6480 -88405 -6392
rect -86235 -6480 -86095 -6290
rect -84015 -6392 -83995 -2248
rect -83895 -6392 -83875 -2248
rect -81705 -2350 -81565 -1970
rect -79485 -2072 -79465 2072
rect -79365 -2072 -79345 2072
rect -77175 1970 -77035 2350
rect -74955 2248 -74935 6392
rect -74835 2248 -74815 6392
rect -72645 6290 -72505 6480
rect -70425 6392 -70285 6480
rect -74955 2072 -74815 2248
rect -79485 -2248 -79345 -2072
rect -84015 -6480 -83875 -6392
rect -81705 -6480 -81565 -6290
rect -79485 -6392 -79465 -2248
rect -79365 -6392 -79345 -2248
rect -77175 -2350 -77035 -1970
rect -74955 -2072 -74935 2072
rect -74835 -2072 -74815 2072
rect -72645 1970 -72505 2350
rect -70425 2248 -70405 6392
rect -70305 2248 -70285 6392
rect -68115 6290 -67975 6480
rect -65895 6392 -65755 6480
rect -70425 2072 -70285 2248
rect -74955 -2248 -74815 -2072
rect -79485 -6480 -79345 -6392
rect -77175 -6480 -77035 -6290
rect -74955 -6392 -74935 -2248
rect -74835 -6392 -74815 -2248
rect -72645 -2350 -72505 -1970
rect -70425 -2072 -70405 2072
rect -70305 -2072 -70285 2072
rect -68115 1970 -67975 2350
rect -65895 2248 -65875 6392
rect -65775 2248 -65755 6392
rect -63585 6290 -63445 6480
rect -61365 6392 -61225 6480
rect -65895 2072 -65755 2248
rect -70425 -2248 -70285 -2072
rect -74955 -6480 -74815 -6392
rect -72645 -6480 -72505 -6290
rect -70425 -6392 -70405 -2248
rect -70305 -6392 -70285 -2248
rect -68115 -2350 -67975 -1970
rect -65895 -2072 -65875 2072
rect -65775 -2072 -65755 2072
rect -63585 1970 -63445 2350
rect -61365 2248 -61345 6392
rect -61245 2248 -61225 6392
rect -59055 6290 -58915 6480
rect -56835 6392 -56695 6480
rect -61365 2072 -61225 2248
rect -65895 -2248 -65755 -2072
rect -70425 -6480 -70285 -6392
rect -68115 -6480 -67975 -6290
rect -65895 -6392 -65875 -2248
rect -65775 -6392 -65755 -2248
rect -63585 -2350 -63445 -1970
rect -61365 -2072 -61345 2072
rect -61245 -2072 -61225 2072
rect -59055 1970 -58915 2350
rect -56835 2248 -56815 6392
rect -56715 2248 -56695 6392
rect -54525 6290 -54385 6480
rect -52305 6392 -52165 6480
rect -56835 2072 -56695 2248
rect -61365 -2248 -61225 -2072
rect -65895 -6480 -65755 -6392
rect -63585 -6480 -63445 -6290
rect -61365 -6392 -61345 -2248
rect -61245 -6392 -61225 -2248
rect -59055 -2350 -58915 -1970
rect -56835 -2072 -56815 2072
rect -56715 -2072 -56695 2072
rect -54525 1970 -54385 2350
rect -52305 2248 -52285 6392
rect -52185 2248 -52165 6392
rect -49995 6290 -49855 6480
rect -47775 6392 -47635 6480
rect -52305 2072 -52165 2248
rect -56835 -2248 -56695 -2072
rect -61365 -6480 -61225 -6392
rect -59055 -6480 -58915 -6290
rect -56835 -6392 -56815 -2248
rect -56715 -6392 -56695 -2248
rect -54525 -2350 -54385 -1970
rect -52305 -2072 -52285 2072
rect -52185 -2072 -52165 2072
rect -49995 1970 -49855 2350
rect -47775 2248 -47755 6392
rect -47655 2248 -47635 6392
rect -45465 6290 -45325 6480
rect -43245 6392 -43105 6480
rect -47775 2072 -47635 2248
rect -52305 -2248 -52165 -2072
rect -56835 -6480 -56695 -6392
rect -54525 -6480 -54385 -6290
rect -52305 -6392 -52285 -2248
rect -52185 -6392 -52165 -2248
rect -49995 -2350 -49855 -1970
rect -47775 -2072 -47755 2072
rect -47655 -2072 -47635 2072
rect -45465 1970 -45325 2350
rect -43245 2248 -43225 6392
rect -43125 2248 -43105 6392
rect -40935 6290 -40795 6480
rect -38715 6392 -38575 6480
rect -43245 2072 -43105 2248
rect -47775 -2248 -47635 -2072
rect -52305 -6480 -52165 -6392
rect -49995 -6480 -49855 -6290
rect -47775 -6392 -47755 -2248
rect -47655 -6392 -47635 -2248
rect -45465 -2350 -45325 -1970
rect -43245 -2072 -43225 2072
rect -43125 -2072 -43105 2072
rect -40935 1970 -40795 2350
rect -38715 2248 -38695 6392
rect -38595 2248 -38575 6392
rect -36405 6290 -36265 6480
rect -34185 6392 -34045 6480
rect -38715 2072 -38575 2248
rect -43245 -2248 -43105 -2072
rect -47775 -6480 -47635 -6392
rect -45465 -6480 -45325 -6290
rect -43245 -6392 -43225 -2248
rect -43125 -6392 -43105 -2248
rect -40935 -2350 -40795 -1970
rect -38715 -2072 -38695 2072
rect -38595 -2072 -38575 2072
rect -36405 1970 -36265 2350
rect -34185 2248 -34165 6392
rect -34065 2248 -34045 6392
rect -31875 6290 -31735 6480
rect -29655 6392 -29515 6480
rect -34185 2072 -34045 2248
rect -38715 -2248 -38575 -2072
rect -43245 -6480 -43105 -6392
rect -40935 -6480 -40795 -6290
rect -38715 -6392 -38695 -2248
rect -38595 -6392 -38575 -2248
rect -36405 -2350 -36265 -1970
rect -34185 -2072 -34165 2072
rect -34065 -2072 -34045 2072
rect -31875 1970 -31735 2350
rect -29655 2248 -29635 6392
rect -29535 2248 -29515 6392
rect -27345 6290 -27205 6480
rect -25125 6392 -24985 6480
rect -29655 2072 -29515 2248
rect -34185 -2248 -34045 -2072
rect -38715 -6480 -38575 -6392
rect -36405 -6480 -36265 -6290
rect -34185 -6392 -34165 -2248
rect -34065 -6392 -34045 -2248
rect -31875 -2350 -31735 -1970
rect -29655 -2072 -29635 2072
rect -29535 -2072 -29515 2072
rect -27345 1970 -27205 2350
rect -25125 2248 -25105 6392
rect -25005 2248 -24985 6392
rect -22815 6290 -22675 6480
rect -20595 6392 -20455 6480
rect -25125 2072 -24985 2248
rect -29655 -2248 -29515 -2072
rect -34185 -6480 -34045 -6392
rect -31875 -6480 -31735 -6290
rect -29655 -6392 -29635 -2248
rect -29535 -6392 -29515 -2248
rect -27345 -2350 -27205 -1970
rect -25125 -2072 -25105 2072
rect -25005 -2072 -24985 2072
rect -22815 1970 -22675 2350
rect -20595 2248 -20575 6392
rect -20475 2248 -20455 6392
rect -18285 6290 -18145 6480
rect -16065 6392 -15925 6480
rect -20595 2072 -20455 2248
rect -25125 -2248 -24985 -2072
rect -29655 -6480 -29515 -6392
rect -27345 -6480 -27205 -6290
rect -25125 -6392 -25105 -2248
rect -25005 -6392 -24985 -2248
rect -22815 -2350 -22675 -1970
rect -20595 -2072 -20575 2072
rect -20475 -2072 -20455 2072
rect -18285 1970 -18145 2350
rect -16065 2248 -16045 6392
rect -15945 2248 -15925 6392
rect -13755 6290 -13615 6480
rect -11535 6392 -11395 6480
rect -16065 2072 -15925 2248
rect -20595 -2248 -20455 -2072
rect -25125 -6480 -24985 -6392
rect -22815 -6480 -22675 -6290
rect -20595 -6392 -20575 -2248
rect -20475 -6392 -20455 -2248
rect -18285 -2350 -18145 -1970
rect -16065 -2072 -16045 2072
rect -15945 -2072 -15925 2072
rect -13755 1970 -13615 2350
rect -11535 2248 -11515 6392
rect -11415 2248 -11395 6392
rect -9225 6290 -9085 6480
rect -7005 6392 -6865 6480
rect -11535 2072 -11395 2248
rect -16065 -2248 -15925 -2072
rect -20595 -6480 -20455 -6392
rect -18285 -6480 -18145 -6290
rect -16065 -6392 -16045 -2248
rect -15945 -6392 -15925 -2248
rect -13755 -2350 -13615 -1970
rect -11535 -2072 -11515 2072
rect -11415 -2072 -11395 2072
rect -9225 1970 -9085 2350
rect -7005 2248 -6985 6392
rect -6885 2248 -6865 6392
rect -4695 6290 -4555 6480
rect -2475 6392 -2335 6480
rect -7005 2072 -6865 2248
rect -11535 -2248 -11395 -2072
rect -16065 -6480 -15925 -6392
rect -13755 -6480 -13615 -6290
rect -11535 -6392 -11515 -2248
rect -11415 -6392 -11395 -2248
rect -9225 -2350 -9085 -1970
rect -7005 -2072 -6985 2072
rect -6885 -2072 -6865 2072
rect -4695 1970 -4555 2350
rect -2475 2248 -2455 6392
rect -2355 2248 -2335 6392
rect -165 6290 -25 6480
rect 2055 6392 2195 6480
rect -2475 2072 -2335 2248
rect -7005 -2248 -6865 -2072
rect -11535 -6480 -11395 -6392
rect -9225 -6480 -9085 -6290
rect -7005 -6392 -6985 -2248
rect -6885 -6392 -6865 -2248
rect -4695 -2350 -4555 -1970
rect -2475 -2072 -2455 2072
rect -2355 -2072 -2335 2072
rect -165 1970 -25 2350
rect 2055 2248 2075 6392
rect 2175 2248 2195 6392
rect 4365 6290 4505 6480
rect 6585 6392 6725 6480
rect 2055 2072 2195 2248
rect -2475 -2248 -2335 -2072
rect -7005 -6480 -6865 -6392
rect -4695 -6480 -4555 -6290
rect -2475 -6392 -2455 -2248
rect -2355 -6392 -2335 -2248
rect -165 -2350 -25 -1970
rect 2055 -2072 2075 2072
rect 2175 -2072 2195 2072
rect 4365 1970 4505 2350
rect 6585 2248 6605 6392
rect 6705 2248 6725 6392
rect 8895 6290 9035 6480
rect 11115 6392 11255 6480
rect 6585 2072 6725 2248
rect 2055 -2248 2195 -2072
rect -2475 -6480 -2335 -6392
rect -165 -6480 -25 -6290
rect 2055 -6392 2075 -2248
rect 2175 -6392 2195 -2248
rect 4365 -2350 4505 -1970
rect 6585 -2072 6605 2072
rect 6705 -2072 6725 2072
rect 8895 1970 9035 2350
rect 11115 2248 11135 6392
rect 11235 2248 11255 6392
rect 13425 6290 13565 6480
rect 15645 6392 15785 6480
rect 11115 2072 11255 2248
rect 6585 -2248 6725 -2072
rect 2055 -6480 2195 -6392
rect 4365 -6480 4505 -6290
rect 6585 -6392 6605 -2248
rect 6705 -6392 6725 -2248
rect 8895 -2350 9035 -1970
rect 11115 -2072 11135 2072
rect 11235 -2072 11255 2072
rect 13425 1970 13565 2350
rect 15645 2248 15665 6392
rect 15765 2248 15785 6392
rect 17955 6290 18095 6480
rect 20175 6392 20315 6480
rect 15645 2072 15785 2248
rect 11115 -2248 11255 -2072
rect 6585 -6480 6725 -6392
rect 8895 -6480 9035 -6290
rect 11115 -6392 11135 -2248
rect 11235 -6392 11255 -2248
rect 13425 -2350 13565 -1970
rect 15645 -2072 15665 2072
rect 15765 -2072 15785 2072
rect 17955 1970 18095 2350
rect 20175 2248 20195 6392
rect 20295 2248 20315 6392
rect 22485 6290 22625 6480
rect 24705 6392 24845 6480
rect 20175 2072 20315 2248
rect 15645 -2248 15785 -2072
rect 11115 -6480 11255 -6392
rect 13425 -6480 13565 -6290
rect 15645 -6392 15665 -2248
rect 15765 -6392 15785 -2248
rect 17955 -2350 18095 -1970
rect 20175 -2072 20195 2072
rect 20295 -2072 20315 2072
rect 22485 1970 22625 2350
rect 24705 2248 24725 6392
rect 24825 2248 24845 6392
rect 27015 6290 27155 6480
rect 29235 6392 29375 6480
rect 24705 2072 24845 2248
rect 20175 -2248 20315 -2072
rect 15645 -6480 15785 -6392
rect 17955 -6480 18095 -6290
rect 20175 -6392 20195 -2248
rect 20295 -6392 20315 -2248
rect 22485 -2350 22625 -1970
rect 24705 -2072 24725 2072
rect 24825 -2072 24845 2072
rect 27015 1970 27155 2350
rect 29235 2248 29255 6392
rect 29355 2248 29375 6392
rect 31545 6290 31685 6480
rect 33765 6392 33905 6480
rect 29235 2072 29375 2248
rect 24705 -2248 24845 -2072
rect 20175 -6480 20315 -6392
rect 22485 -6480 22625 -6290
rect 24705 -6392 24725 -2248
rect 24825 -6392 24845 -2248
rect 27015 -2350 27155 -1970
rect 29235 -2072 29255 2072
rect 29355 -2072 29375 2072
rect 31545 1970 31685 2350
rect 33765 2248 33785 6392
rect 33885 2248 33905 6392
rect 36075 6290 36215 6480
rect 38295 6392 38435 6480
rect 33765 2072 33905 2248
rect 29235 -2248 29375 -2072
rect 24705 -6480 24845 -6392
rect 27015 -6480 27155 -6290
rect 29235 -6392 29255 -2248
rect 29355 -6392 29375 -2248
rect 31545 -2350 31685 -1970
rect 33765 -2072 33785 2072
rect 33885 -2072 33905 2072
rect 36075 1970 36215 2350
rect 38295 2248 38315 6392
rect 38415 2248 38435 6392
rect 40605 6290 40745 6480
rect 42825 6392 42965 6480
rect 38295 2072 38435 2248
rect 33765 -2248 33905 -2072
rect 29235 -6480 29375 -6392
rect 31545 -6480 31685 -6290
rect 33765 -6392 33785 -2248
rect 33885 -6392 33905 -2248
rect 36075 -2350 36215 -1970
rect 38295 -2072 38315 2072
rect 38415 -2072 38435 2072
rect 40605 1970 40745 2350
rect 42825 2248 42845 6392
rect 42945 2248 42965 6392
rect 45135 6290 45275 6480
rect 47355 6392 47495 6480
rect 42825 2072 42965 2248
rect 38295 -2248 38435 -2072
rect 33765 -6480 33905 -6392
rect 36075 -6480 36215 -6290
rect 38295 -6392 38315 -2248
rect 38415 -6392 38435 -2248
rect 40605 -2350 40745 -1970
rect 42825 -2072 42845 2072
rect 42945 -2072 42965 2072
rect 45135 1970 45275 2350
rect 47355 2248 47375 6392
rect 47475 2248 47495 6392
rect 49665 6290 49805 6480
rect 51885 6392 52025 6480
rect 47355 2072 47495 2248
rect 42825 -2248 42965 -2072
rect 38295 -6480 38435 -6392
rect 40605 -6480 40745 -6290
rect 42825 -6392 42845 -2248
rect 42945 -6392 42965 -2248
rect 45135 -2350 45275 -1970
rect 47355 -2072 47375 2072
rect 47475 -2072 47495 2072
rect 49665 1970 49805 2350
rect 51885 2248 51905 6392
rect 52005 2248 52025 6392
rect 54195 6290 54335 6480
rect 56415 6392 56555 6480
rect 51885 2072 52025 2248
rect 47355 -2248 47495 -2072
rect 42825 -6480 42965 -6392
rect 45135 -6480 45275 -6290
rect 47355 -6392 47375 -2248
rect 47475 -6392 47495 -2248
rect 49665 -2350 49805 -1970
rect 51885 -2072 51905 2072
rect 52005 -2072 52025 2072
rect 54195 1970 54335 2350
rect 56415 2248 56435 6392
rect 56535 2248 56555 6392
rect 58725 6290 58865 6480
rect 60945 6392 61085 6480
rect 56415 2072 56555 2248
rect 51885 -2248 52025 -2072
rect 47355 -6480 47495 -6392
rect 49665 -6480 49805 -6290
rect 51885 -6392 51905 -2248
rect 52005 -6392 52025 -2248
rect 54195 -2350 54335 -1970
rect 56415 -2072 56435 2072
rect 56535 -2072 56555 2072
rect 58725 1970 58865 2350
rect 60945 2248 60965 6392
rect 61065 2248 61085 6392
rect 63255 6290 63395 6480
rect 65475 6392 65615 6480
rect 60945 2072 61085 2248
rect 56415 -2248 56555 -2072
rect 51885 -6480 52025 -6392
rect 54195 -6480 54335 -6290
rect 56415 -6392 56435 -2248
rect 56535 -6392 56555 -2248
rect 58725 -2350 58865 -1970
rect 60945 -2072 60965 2072
rect 61065 -2072 61085 2072
rect 63255 1970 63395 2350
rect 65475 2248 65495 6392
rect 65595 2248 65615 6392
rect 67785 6290 67925 6480
rect 70005 6392 70145 6480
rect 65475 2072 65615 2248
rect 60945 -2248 61085 -2072
rect 56415 -6480 56555 -6392
rect 58725 -6480 58865 -6290
rect 60945 -6392 60965 -2248
rect 61065 -6392 61085 -2248
rect 63255 -2350 63395 -1970
rect 65475 -2072 65495 2072
rect 65595 -2072 65615 2072
rect 67785 1970 67925 2350
rect 70005 2248 70025 6392
rect 70125 2248 70145 6392
rect 72315 6290 72455 6480
rect 74535 6392 74675 6480
rect 70005 2072 70145 2248
rect 65475 -2248 65615 -2072
rect 60945 -6480 61085 -6392
rect 63255 -6480 63395 -6290
rect 65475 -6392 65495 -2248
rect 65595 -6392 65615 -2248
rect 67785 -2350 67925 -1970
rect 70005 -2072 70025 2072
rect 70125 -2072 70145 2072
rect 72315 1970 72455 2350
rect 74535 2248 74555 6392
rect 74655 2248 74675 6392
rect 76845 6290 76985 6480
rect 79065 6392 79205 6480
rect 74535 2072 74675 2248
rect 70005 -2248 70145 -2072
rect 65475 -6480 65615 -6392
rect 67785 -6480 67925 -6290
rect 70005 -6392 70025 -2248
rect 70125 -6392 70145 -2248
rect 72315 -2350 72455 -1970
rect 74535 -2072 74555 2072
rect 74655 -2072 74675 2072
rect 76845 1970 76985 2350
rect 79065 2248 79085 6392
rect 79185 2248 79205 6392
rect 81375 6290 81515 6480
rect 83595 6392 83735 6480
rect 79065 2072 79205 2248
rect 74535 -2248 74675 -2072
rect 70005 -6480 70145 -6392
rect 72315 -6480 72455 -6290
rect 74535 -6392 74555 -2248
rect 74655 -6392 74675 -2248
rect 76845 -2350 76985 -1970
rect 79065 -2072 79085 2072
rect 79185 -2072 79205 2072
rect 81375 1970 81515 2350
rect 83595 2248 83615 6392
rect 83715 2248 83735 6392
rect 85905 6290 86045 6480
rect 88125 6392 88265 6480
rect 83595 2072 83735 2248
rect 79065 -2248 79205 -2072
rect 74535 -6480 74675 -6392
rect 76845 -6480 76985 -6290
rect 79065 -6392 79085 -2248
rect 79185 -6392 79205 -2248
rect 81375 -2350 81515 -1970
rect 83595 -2072 83615 2072
rect 83715 -2072 83735 2072
rect 85905 1970 86045 2350
rect 88125 2248 88145 6392
rect 88245 2248 88265 6392
rect 90435 6290 90575 6480
rect 92655 6392 92795 6480
rect 88125 2072 88265 2248
rect 83595 -2248 83735 -2072
rect 79065 -6480 79205 -6392
rect 81375 -6480 81515 -6290
rect 83595 -6392 83615 -2248
rect 83715 -6392 83735 -2248
rect 85905 -2350 86045 -1970
rect 88125 -2072 88145 2072
rect 88245 -2072 88265 2072
rect 90435 1970 90575 2350
rect 92655 2248 92675 6392
rect 92775 2248 92795 6392
rect 94965 6290 95105 6480
rect 97185 6392 97325 6480
rect 92655 2072 92795 2248
rect 88125 -2248 88265 -2072
rect 83595 -6480 83735 -6392
rect 85905 -6480 86045 -6290
rect 88125 -6392 88145 -2248
rect 88245 -6392 88265 -2248
rect 90435 -2350 90575 -1970
rect 92655 -2072 92675 2072
rect 92775 -2072 92795 2072
rect 94965 1970 95105 2350
rect 97185 2248 97205 6392
rect 97305 2248 97325 6392
rect 99495 6290 99635 6480
rect 101715 6392 101855 6480
rect 97185 2072 97325 2248
rect 92655 -2248 92795 -2072
rect 88125 -6480 88265 -6392
rect 90435 -6480 90575 -6290
rect 92655 -6392 92675 -2248
rect 92775 -6392 92795 -2248
rect 94965 -2350 95105 -1970
rect 97185 -2072 97205 2072
rect 97305 -2072 97325 2072
rect 99495 1970 99635 2350
rect 101715 2248 101735 6392
rect 101835 2248 101855 6392
rect 104025 6290 104165 6480
rect 106245 6392 106385 6480
rect 101715 2072 101855 2248
rect 97185 -2248 97325 -2072
rect 92655 -6480 92795 -6392
rect 94965 -6480 95105 -6290
rect 97185 -6392 97205 -2248
rect 97305 -6392 97325 -2248
rect 99495 -2350 99635 -1970
rect 101715 -2072 101735 2072
rect 101835 -2072 101855 2072
rect 104025 1970 104165 2350
rect 106245 2248 106265 6392
rect 106365 2248 106385 6392
rect 108555 6290 108695 6480
rect 110775 6392 110915 6480
rect 106245 2072 106385 2248
rect 101715 -2248 101855 -2072
rect 97185 -6480 97325 -6392
rect 99495 -6480 99635 -6290
rect 101715 -6392 101735 -2248
rect 101835 -6392 101855 -2248
rect 104025 -2350 104165 -1970
rect 106245 -2072 106265 2072
rect 106365 -2072 106385 2072
rect 108555 1970 108695 2350
rect 110775 2248 110795 6392
rect 110895 2248 110915 6392
rect 113085 6290 113225 6480
rect 115305 6392 115445 6480
rect 110775 2072 110915 2248
rect 106245 -2248 106385 -2072
rect 101715 -6480 101855 -6392
rect 104025 -6480 104165 -6290
rect 106245 -6392 106265 -2248
rect 106365 -6392 106385 -2248
rect 108555 -2350 108695 -1970
rect 110775 -2072 110795 2072
rect 110895 -2072 110915 2072
rect 113085 1970 113225 2350
rect 115305 2248 115325 6392
rect 115425 2248 115445 6392
rect 117615 6290 117755 6480
rect 119835 6392 119975 6480
rect 115305 2072 115445 2248
rect 110775 -2248 110915 -2072
rect 106245 -6480 106385 -6392
rect 108555 -6480 108695 -6290
rect 110775 -6392 110795 -2248
rect 110895 -6392 110915 -2248
rect 113085 -2350 113225 -1970
rect 115305 -2072 115325 2072
rect 115425 -2072 115445 2072
rect 117615 1970 117755 2350
rect 119835 2248 119855 6392
rect 119955 2248 119975 6392
rect 122145 6290 122285 6480
rect 124365 6392 124505 6480
rect 119835 2072 119975 2248
rect 115305 -2248 115445 -2072
rect 110775 -6480 110915 -6392
rect 113085 -6480 113225 -6290
rect 115305 -6392 115325 -2248
rect 115425 -6392 115445 -2248
rect 117615 -2350 117755 -1970
rect 119835 -2072 119855 2072
rect 119955 -2072 119975 2072
rect 122145 1970 122285 2350
rect 124365 2248 124385 6392
rect 124485 2248 124505 6392
rect 124365 2072 124505 2248
rect 119835 -2248 119975 -2072
rect 115305 -6480 115445 -6392
rect 117615 -6480 117755 -6290
rect 119835 -6392 119855 -2248
rect 119955 -6392 119975 -2248
rect 122145 -2350 122285 -1970
rect 124365 -2072 124385 2072
rect 124485 -2072 124505 2072
rect 124365 -2248 124505 -2072
rect 119835 -6480 119975 -6392
rect 122145 -6480 122285 -6290
rect 124365 -6392 124385 -2248
rect 124485 -6392 124505 -2248
rect 124365 -6480 124505 -6392
<< properties >>
string parameters w 20.00 l 20.00 val 413.6 carea 1.00 cperi 0.17 nx 55 ny 3 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
