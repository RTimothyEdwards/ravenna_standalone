magic
tech EFXH018D
timestamp 1494891594
<< metal2 >>
rect 0 848 528 960
rect 0 528 96 848
rect 0 416 368 528
rect 0 0 96 416
<< end >>
