magic
tech EFXH018D
timestamp 1565723183
<< mimcap >>
rect -2180 60385 -180 60400
rect -2180 58415 -2165 60385
rect -195 58415 -180 60385
rect -2180 58400 -180 58415
rect 85 60385 2085 60400
rect 85 58415 100 60385
rect 2070 58415 2085 60385
rect 85 58400 2085 58415
rect -2180 58225 -180 58240
rect -2180 56255 -2165 58225
rect -195 56255 -180 58225
rect -2180 56240 -180 56255
rect 85 58225 2085 58240
rect 85 56255 100 58225
rect 2070 56255 2085 58225
rect 85 56240 2085 56255
rect -2180 56065 -180 56080
rect -2180 54095 -2165 56065
rect -195 54095 -180 56065
rect -2180 54080 -180 54095
rect 85 56065 2085 56080
rect 85 54095 100 56065
rect 2070 54095 2085 56065
rect 85 54080 2085 54095
rect -2180 53905 -180 53920
rect -2180 51935 -2165 53905
rect -195 51935 -180 53905
rect -2180 51920 -180 51935
rect 85 53905 2085 53920
rect 85 51935 100 53905
rect 2070 51935 2085 53905
rect 85 51920 2085 51935
rect -2180 51745 -180 51760
rect -2180 49775 -2165 51745
rect -195 49775 -180 51745
rect -2180 49760 -180 49775
rect 85 51745 2085 51760
rect 85 49775 100 51745
rect 2070 49775 2085 51745
rect 85 49760 2085 49775
rect -2180 49585 -180 49600
rect -2180 47615 -2165 49585
rect -195 47615 -180 49585
rect -2180 47600 -180 47615
rect 85 49585 2085 49600
rect 85 47615 100 49585
rect 2070 47615 2085 49585
rect 85 47600 2085 47615
rect -2180 47425 -180 47440
rect -2180 45455 -2165 47425
rect -195 45455 -180 47425
rect -2180 45440 -180 45455
rect 85 47425 2085 47440
rect 85 45455 100 47425
rect 2070 45455 2085 47425
rect 85 45440 2085 45455
rect -2180 45265 -180 45280
rect -2180 43295 -2165 45265
rect -195 43295 -180 45265
rect -2180 43280 -180 43295
rect 85 45265 2085 45280
rect 85 43295 100 45265
rect 2070 43295 2085 45265
rect 85 43280 2085 43295
rect -2180 43105 -180 43120
rect -2180 41135 -2165 43105
rect -195 41135 -180 43105
rect -2180 41120 -180 41135
rect 85 43105 2085 43120
rect 85 41135 100 43105
rect 2070 41135 2085 43105
rect 85 41120 2085 41135
rect -2180 40945 -180 40960
rect -2180 38975 -2165 40945
rect -195 38975 -180 40945
rect -2180 38960 -180 38975
rect 85 40945 2085 40960
rect 85 38975 100 40945
rect 2070 38975 2085 40945
rect 85 38960 2085 38975
rect -2180 38785 -180 38800
rect -2180 36815 -2165 38785
rect -195 36815 -180 38785
rect -2180 36800 -180 36815
rect 85 38785 2085 38800
rect 85 36815 100 38785
rect 2070 36815 2085 38785
rect 85 36800 2085 36815
rect -2180 36625 -180 36640
rect -2180 34655 -2165 36625
rect -195 34655 -180 36625
rect -2180 34640 -180 34655
rect 85 36625 2085 36640
rect 85 34655 100 36625
rect 2070 34655 2085 36625
rect 85 34640 2085 34655
rect -2180 34465 -180 34480
rect -2180 32495 -2165 34465
rect -195 32495 -180 34465
rect -2180 32480 -180 32495
rect 85 34465 2085 34480
rect 85 32495 100 34465
rect 2070 32495 2085 34465
rect 85 32480 2085 32495
rect -2180 32305 -180 32320
rect -2180 30335 -2165 32305
rect -195 30335 -180 32305
rect -2180 30320 -180 30335
rect 85 32305 2085 32320
rect 85 30335 100 32305
rect 2070 30335 2085 32305
rect 85 30320 2085 30335
rect -2180 30145 -180 30160
rect -2180 28175 -2165 30145
rect -195 28175 -180 30145
rect -2180 28160 -180 28175
rect 85 30145 2085 30160
rect 85 28175 100 30145
rect 2070 28175 2085 30145
rect 85 28160 2085 28175
rect -2180 27985 -180 28000
rect -2180 26015 -2165 27985
rect -195 26015 -180 27985
rect -2180 26000 -180 26015
rect 85 27985 2085 28000
rect 85 26015 100 27985
rect 2070 26015 2085 27985
rect 85 26000 2085 26015
rect -2180 25825 -180 25840
rect -2180 23855 -2165 25825
rect -195 23855 -180 25825
rect -2180 23840 -180 23855
rect 85 25825 2085 25840
rect 85 23855 100 25825
rect 2070 23855 2085 25825
rect 85 23840 2085 23855
rect -2180 23665 -180 23680
rect -2180 21695 -2165 23665
rect -195 21695 -180 23665
rect -2180 21680 -180 21695
rect 85 23665 2085 23680
rect 85 21695 100 23665
rect 2070 21695 2085 23665
rect 85 21680 2085 21695
rect -2180 21505 -180 21520
rect -2180 19535 -2165 21505
rect -195 19535 -180 21505
rect -2180 19520 -180 19535
rect 85 21505 2085 21520
rect 85 19535 100 21505
rect 2070 19535 2085 21505
rect 85 19520 2085 19535
rect -2180 19345 -180 19360
rect -2180 17375 -2165 19345
rect -195 17375 -180 19345
rect -2180 17360 -180 17375
rect 85 19345 2085 19360
rect 85 17375 100 19345
rect 2070 17375 2085 19345
rect 85 17360 2085 17375
rect -2180 17185 -180 17200
rect -2180 15215 -2165 17185
rect -195 15215 -180 17185
rect -2180 15200 -180 15215
rect 85 17185 2085 17200
rect 85 15215 100 17185
rect 2070 15215 2085 17185
rect 85 15200 2085 15215
rect -2180 15025 -180 15040
rect -2180 13055 -2165 15025
rect -195 13055 -180 15025
rect -2180 13040 -180 13055
rect 85 15025 2085 15040
rect 85 13055 100 15025
rect 2070 13055 2085 15025
rect 85 13040 2085 13055
rect -2180 12865 -180 12880
rect -2180 10895 -2165 12865
rect -195 10895 -180 12865
rect -2180 10880 -180 10895
rect 85 12865 2085 12880
rect 85 10895 100 12865
rect 2070 10895 2085 12865
rect 85 10880 2085 10895
rect -2180 10705 -180 10720
rect -2180 8735 -2165 10705
rect -195 8735 -180 10705
rect -2180 8720 -180 8735
rect 85 10705 2085 10720
rect 85 8735 100 10705
rect 2070 8735 2085 10705
rect 85 8720 2085 8735
rect -2180 8545 -180 8560
rect -2180 6575 -2165 8545
rect -195 6575 -180 8545
rect -2180 6560 -180 6575
rect 85 8545 2085 8560
rect 85 6575 100 8545
rect 2070 6575 2085 8545
rect 85 6560 2085 6575
rect -2180 6385 -180 6400
rect -2180 4415 -2165 6385
rect -195 4415 -180 6385
rect -2180 4400 -180 4415
rect 85 6385 2085 6400
rect 85 4415 100 6385
rect 2070 4415 2085 6385
rect 85 4400 2085 4415
rect -2180 4225 -180 4240
rect -2180 2255 -2165 4225
rect -195 2255 -180 4225
rect -2180 2240 -180 2255
rect 85 4225 2085 4240
rect 85 2255 100 4225
rect 2070 2255 2085 4225
rect 85 2240 2085 2255
rect -2180 2065 -180 2080
rect -2180 95 -2165 2065
rect -195 95 -180 2065
rect -2180 80 -180 95
rect 85 2065 2085 2080
rect 85 95 100 2065
rect 2070 95 2085 2065
rect 85 80 2085 95
rect -2180 -95 -180 -80
rect -2180 -2065 -2165 -95
rect -195 -2065 -180 -95
rect -2180 -2080 -180 -2065
rect 85 -95 2085 -80
rect 85 -2065 100 -95
rect 2070 -2065 2085 -95
rect 85 -2080 2085 -2065
rect -2180 -2255 -180 -2240
rect -2180 -4225 -2165 -2255
rect -195 -4225 -180 -2255
rect -2180 -4240 -180 -4225
rect 85 -2255 2085 -2240
rect 85 -4225 100 -2255
rect 2070 -4225 2085 -2255
rect 85 -4240 2085 -4225
rect -2180 -4415 -180 -4400
rect -2180 -6385 -2165 -4415
rect -195 -6385 -180 -4415
rect -2180 -6400 -180 -6385
rect 85 -4415 2085 -4400
rect 85 -6385 100 -4415
rect 2070 -6385 2085 -4415
rect 85 -6400 2085 -6385
rect -2180 -6575 -180 -6560
rect -2180 -8545 -2165 -6575
rect -195 -8545 -180 -6575
rect -2180 -8560 -180 -8545
rect 85 -6575 2085 -6560
rect 85 -8545 100 -6575
rect 2070 -8545 2085 -6575
rect 85 -8560 2085 -8545
rect -2180 -8735 -180 -8720
rect -2180 -10705 -2165 -8735
rect -195 -10705 -180 -8735
rect -2180 -10720 -180 -10705
rect 85 -8735 2085 -8720
rect 85 -10705 100 -8735
rect 2070 -10705 2085 -8735
rect 85 -10720 2085 -10705
rect -2180 -10895 -180 -10880
rect -2180 -12865 -2165 -10895
rect -195 -12865 -180 -10895
rect -2180 -12880 -180 -12865
rect 85 -10895 2085 -10880
rect 85 -12865 100 -10895
rect 2070 -12865 2085 -10895
rect 85 -12880 2085 -12865
rect -2180 -13055 -180 -13040
rect -2180 -15025 -2165 -13055
rect -195 -15025 -180 -13055
rect -2180 -15040 -180 -15025
rect 85 -13055 2085 -13040
rect 85 -15025 100 -13055
rect 2070 -15025 2085 -13055
rect 85 -15040 2085 -15025
rect -2180 -15215 -180 -15200
rect -2180 -17185 -2165 -15215
rect -195 -17185 -180 -15215
rect -2180 -17200 -180 -17185
rect 85 -15215 2085 -15200
rect 85 -17185 100 -15215
rect 2070 -17185 2085 -15215
rect 85 -17200 2085 -17185
rect -2180 -17375 -180 -17360
rect -2180 -19345 -2165 -17375
rect -195 -19345 -180 -17375
rect -2180 -19360 -180 -19345
rect 85 -17375 2085 -17360
rect 85 -19345 100 -17375
rect 2070 -19345 2085 -17375
rect 85 -19360 2085 -19345
rect -2180 -19535 -180 -19520
rect -2180 -21505 -2165 -19535
rect -195 -21505 -180 -19535
rect -2180 -21520 -180 -21505
rect 85 -19535 2085 -19520
rect 85 -21505 100 -19535
rect 2070 -21505 2085 -19535
rect 85 -21520 2085 -21505
rect -2180 -21695 -180 -21680
rect -2180 -23665 -2165 -21695
rect -195 -23665 -180 -21695
rect -2180 -23680 -180 -23665
rect 85 -21695 2085 -21680
rect 85 -23665 100 -21695
rect 2070 -23665 2085 -21695
rect 85 -23680 2085 -23665
rect -2180 -23855 -180 -23840
rect -2180 -25825 -2165 -23855
rect -195 -25825 -180 -23855
rect -2180 -25840 -180 -25825
rect 85 -23855 2085 -23840
rect 85 -25825 100 -23855
rect 2070 -25825 2085 -23855
rect 85 -25840 2085 -25825
rect -2180 -26015 -180 -26000
rect -2180 -27985 -2165 -26015
rect -195 -27985 -180 -26015
rect -2180 -28000 -180 -27985
rect 85 -26015 2085 -26000
rect 85 -27985 100 -26015
rect 2070 -27985 2085 -26015
rect 85 -28000 2085 -27985
rect -2180 -28175 -180 -28160
rect -2180 -30145 -2165 -28175
rect -195 -30145 -180 -28175
rect -2180 -30160 -180 -30145
rect 85 -28175 2085 -28160
rect 85 -30145 100 -28175
rect 2070 -30145 2085 -28175
rect 85 -30160 2085 -30145
rect -2180 -30335 -180 -30320
rect -2180 -32305 -2165 -30335
rect -195 -32305 -180 -30335
rect -2180 -32320 -180 -32305
rect 85 -30335 2085 -30320
rect 85 -32305 100 -30335
rect 2070 -32305 2085 -30335
rect 85 -32320 2085 -32305
rect -2180 -32495 -180 -32480
rect -2180 -34465 -2165 -32495
rect -195 -34465 -180 -32495
rect -2180 -34480 -180 -34465
rect 85 -32495 2085 -32480
rect 85 -34465 100 -32495
rect 2070 -34465 2085 -32495
rect 85 -34480 2085 -34465
rect -2180 -34655 -180 -34640
rect -2180 -36625 -2165 -34655
rect -195 -36625 -180 -34655
rect -2180 -36640 -180 -36625
rect 85 -34655 2085 -34640
rect 85 -36625 100 -34655
rect 2070 -36625 2085 -34655
rect 85 -36640 2085 -36625
rect -2180 -36815 -180 -36800
rect -2180 -38785 -2165 -36815
rect -195 -38785 -180 -36815
rect -2180 -38800 -180 -38785
rect 85 -36815 2085 -36800
rect 85 -38785 100 -36815
rect 2070 -38785 2085 -36815
rect 85 -38800 2085 -38785
rect -2180 -38975 -180 -38960
rect -2180 -40945 -2165 -38975
rect -195 -40945 -180 -38975
rect -2180 -40960 -180 -40945
rect 85 -38975 2085 -38960
rect 85 -40945 100 -38975
rect 2070 -40945 2085 -38975
rect 85 -40960 2085 -40945
rect -2180 -41135 -180 -41120
rect -2180 -43105 -2165 -41135
rect -195 -43105 -180 -41135
rect -2180 -43120 -180 -43105
rect 85 -41135 2085 -41120
rect 85 -43105 100 -41135
rect 2070 -43105 2085 -41135
rect 85 -43120 2085 -43105
rect -2180 -43295 -180 -43280
rect -2180 -45265 -2165 -43295
rect -195 -45265 -180 -43295
rect -2180 -45280 -180 -45265
rect 85 -43295 2085 -43280
rect 85 -45265 100 -43295
rect 2070 -45265 2085 -43295
rect 85 -45280 2085 -45265
rect -2180 -45455 -180 -45440
rect -2180 -47425 -2165 -45455
rect -195 -47425 -180 -45455
rect -2180 -47440 -180 -47425
rect 85 -45455 2085 -45440
rect 85 -47425 100 -45455
rect 2070 -47425 2085 -45455
rect 85 -47440 2085 -47425
rect -2180 -47615 -180 -47600
rect -2180 -49585 -2165 -47615
rect -195 -49585 -180 -47615
rect -2180 -49600 -180 -49585
rect 85 -47615 2085 -47600
rect 85 -49585 100 -47615
rect 2070 -49585 2085 -47615
rect 85 -49600 2085 -49585
rect -2180 -49775 -180 -49760
rect -2180 -51745 -2165 -49775
rect -195 -51745 -180 -49775
rect -2180 -51760 -180 -51745
rect 85 -49775 2085 -49760
rect 85 -51745 100 -49775
rect 2070 -51745 2085 -49775
rect 85 -51760 2085 -51745
rect -2180 -51935 -180 -51920
rect -2180 -53905 -2165 -51935
rect -195 -53905 -180 -51935
rect -2180 -53920 -180 -53905
rect 85 -51935 2085 -51920
rect 85 -53905 100 -51935
rect 2070 -53905 2085 -51935
rect 85 -53920 2085 -53905
rect -2180 -54095 -180 -54080
rect -2180 -56065 -2165 -54095
rect -195 -56065 -180 -54095
rect -2180 -56080 -180 -56065
rect 85 -54095 2085 -54080
rect 85 -56065 100 -54095
rect 2070 -56065 2085 -54095
rect 85 -56080 2085 -56065
rect -2180 -56255 -180 -56240
rect -2180 -58225 -2165 -56255
rect -195 -58225 -180 -56255
rect -2180 -58240 -180 -58225
rect 85 -56255 2085 -56240
rect 85 -58225 100 -56255
rect 2070 -58225 2085 -56255
rect 85 -58240 2085 -58225
rect -2180 -58415 -180 -58400
rect -2180 -60385 -2165 -58415
rect -195 -60385 -180 -58415
rect -2180 -60400 -180 -60385
rect 85 -58415 2085 -58400
rect 85 -60385 100 -58415
rect 2070 -60385 2085 -58415
rect 85 -60400 2085 -60385
<< mimcapcontact >>
rect -2165 58415 -195 60385
rect 100 58415 2070 60385
rect -2165 56255 -195 58225
rect 100 56255 2070 58225
rect -2165 54095 -195 56065
rect 100 54095 2070 56065
rect -2165 51935 -195 53905
rect 100 51935 2070 53905
rect -2165 49775 -195 51745
rect 100 49775 2070 51745
rect -2165 47615 -195 49585
rect 100 47615 2070 49585
rect -2165 45455 -195 47425
rect 100 45455 2070 47425
rect -2165 43295 -195 45265
rect 100 43295 2070 45265
rect -2165 41135 -195 43105
rect 100 41135 2070 43105
rect -2165 38975 -195 40945
rect 100 38975 2070 40945
rect -2165 36815 -195 38785
rect 100 36815 2070 38785
rect -2165 34655 -195 36625
rect 100 34655 2070 36625
rect -2165 32495 -195 34465
rect 100 32495 2070 34465
rect -2165 30335 -195 32305
rect 100 30335 2070 32305
rect -2165 28175 -195 30145
rect 100 28175 2070 30145
rect -2165 26015 -195 27985
rect 100 26015 2070 27985
rect -2165 23855 -195 25825
rect 100 23855 2070 25825
rect -2165 21695 -195 23665
rect 100 21695 2070 23665
rect -2165 19535 -195 21505
rect 100 19535 2070 21505
rect -2165 17375 -195 19345
rect 100 17375 2070 19345
rect -2165 15215 -195 17185
rect 100 15215 2070 17185
rect -2165 13055 -195 15025
rect 100 13055 2070 15025
rect -2165 10895 -195 12865
rect 100 10895 2070 12865
rect -2165 8735 -195 10705
rect 100 8735 2070 10705
rect -2165 6575 -195 8545
rect 100 6575 2070 8545
rect -2165 4415 -195 6385
rect 100 4415 2070 6385
rect -2165 2255 -195 4225
rect 100 2255 2070 4225
rect -2165 95 -195 2065
rect 100 95 2070 2065
rect -2165 -2065 -195 -95
rect 100 -2065 2070 -95
rect -2165 -4225 -195 -2255
rect 100 -4225 2070 -2255
rect -2165 -6385 -195 -4415
rect 100 -6385 2070 -4415
rect -2165 -8545 -195 -6575
rect 100 -8545 2070 -6575
rect -2165 -10705 -195 -8735
rect 100 -10705 2070 -8735
rect -2165 -12865 -195 -10895
rect 100 -12865 2070 -10895
rect -2165 -15025 -195 -13055
rect 100 -15025 2070 -13055
rect -2165 -17185 -195 -15215
rect 100 -17185 2070 -15215
rect -2165 -19345 -195 -17375
rect 100 -19345 2070 -17375
rect -2165 -21505 -195 -19535
rect 100 -21505 2070 -19535
rect -2165 -23665 -195 -21695
rect 100 -23665 2070 -21695
rect -2165 -25825 -195 -23855
rect 100 -25825 2070 -23855
rect -2165 -27985 -195 -26015
rect 100 -27985 2070 -26015
rect -2165 -30145 -195 -28175
rect 100 -30145 2070 -28175
rect -2165 -32305 -195 -30335
rect 100 -32305 2070 -30335
rect -2165 -34465 -195 -32495
rect 100 -34465 2070 -32495
rect -2165 -36625 -195 -34655
rect 100 -36625 2070 -34655
rect -2165 -38785 -195 -36815
rect 100 -38785 2070 -36815
rect -2165 -40945 -195 -38975
rect 100 -40945 2070 -38975
rect -2165 -43105 -195 -41135
rect 100 -43105 2070 -41135
rect -2165 -45265 -195 -43295
rect 100 -45265 2070 -43295
rect -2165 -47425 -195 -45455
rect 100 -47425 2070 -45455
rect -2165 -49585 -195 -47615
rect 100 -49585 2070 -47615
rect -2165 -51745 -195 -49775
rect 100 -51745 2070 -49775
rect -2165 -53905 -195 -51935
rect 100 -53905 2070 -51935
rect -2165 -56065 -195 -54095
rect 100 -56065 2070 -54095
rect -2165 -58225 -195 -56255
rect 100 -58225 2070 -56255
rect -2165 -60385 -195 -58415
rect 100 -60385 2070 -58415
<< metal4 >>
rect -2230 60436 -35 60450
rect -2230 60400 -95 60436
rect -2230 58400 -2180 60400
rect -180 58400 -95 60400
rect -2230 58364 -95 58400
rect -45 58364 -35 60436
rect -2230 58350 -35 58364
rect 35 60436 2230 60450
rect 35 60400 2170 60436
rect 35 58400 85 60400
rect 2085 58400 2170 60400
rect 35 58364 2170 58400
rect 2220 58364 2230 60436
rect 35 58350 2230 58364
rect -2230 58276 -35 58290
rect -2230 58240 -95 58276
rect -2230 56240 -2180 58240
rect -180 56240 -95 58240
rect -2230 56204 -95 56240
rect -45 56204 -35 58276
rect -2230 56190 -35 56204
rect 35 58276 2230 58290
rect 35 58240 2170 58276
rect 35 56240 85 58240
rect 2085 56240 2170 58240
rect 35 56204 2170 56240
rect 2220 56204 2230 58276
rect 35 56190 2230 56204
rect -2230 56116 -35 56130
rect -2230 56080 -95 56116
rect -2230 54080 -2180 56080
rect -180 54080 -95 56080
rect -2230 54044 -95 54080
rect -45 54044 -35 56116
rect -2230 54030 -35 54044
rect 35 56116 2230 56130
rect 35 56080 2170 56116
rect 35 54080 85 56080
rect 2085 54080 2170 56080
rect 35 54044 2170 54080
rect 2220 54044 2230 56116
rect 35 54030 2230 54044
rect -2230 53956 -35 53970
rect -2230 53920 -95 53956
rect -2230 51920 -2180 53920
rect -180 51920 -95 53920
rect -2230 51884 -95 51920
rect -45 51884 -35 53956
rect -2230 51870 -35 51884
rect 35 53956 2230 53970
rect 35 53920 2170 53956
rect 35 51920 85 53920
rect 2085 51920 2170 53920
rect 35 51884 2170 51920
rect 2220 51884 2230 53956
rect 35 51870 2230 51884
rect -2230 51796 -35 51810
rect -2230 51760 -95 51796
rect -2230 49760 -2180 51760
rect -180 49760 -95 51760
rect -2230 49724 -95 49760
rect -45 49724 -35 51796
rect -2230 49710 -35 49724
rect 35 51796 2230 51810
rect 35 51760 2170 51796
rect 35 49760 85 51760
rect 2085 49760 2170 51760
rect 35 49724 2170 49760
rect 2220 49724 2230 51796
rect 35 49710 2230 49724
rect -2230 49636 -35 49650
rect -2230 49600 -95 49636
rect -2230 47600 -2180 49600
rect -180 47600 -95 49600
rect -2230 47564 -95 47600
rect -45 47564 -35 49636
rect -2230 47550 -35 47564
rect 35 49636 2230 49650
rect 35 49600 2170 49636
rect 35 47600 85 49600
rect 2085 47600 2170 49600
rect 35 47564 2170 47600
rect 2220 47564 2230 49636
rect 35 47550 2230 47564
rect -2230 47476 -35 47490
rect -2230 47440 -95 47476
rect -2230 45440 -2180 47440
rect -180 45440 -95 47440
rect -2230 45404 -95 45440
rect -45 45404 -35 47476
rect -2230 45390 -35 45404
rect 35 47476 2230 47490
rect 35 47440 2170 47476
rect 35 45440 85 47440
rect 2085 45440 2170 47440
rect 35 45404 2170 45440
rect 2220 45404 2230 47476
rect 35 45390 2230 45404
rect -2230 45316 -35 45330
rect -2230 45280 -95 45316
rect -2230 43280 -2180 45280
rect -180 43280 -95 45280
rect -2230 43244 -95 43280
rect -45 43244 -35 45316
rect -2230 43230 -35 43244
rect 35 45316 2230 45330
rect 35 45280 2170 45316
rect 35 43280 85 45280
rect 2085 43280 2170 45280
rect 35 43244 2170 43280
rect 2220 43244 2230 45316
rect 35 43230 2230 43244
rect -2230 43156 -35 43170
rect -2230 43120 -95 43156
rect -2230 41120 -2180 43120
rect -180 41120 -95 43120
rect -2230 41084 -95 41120
rect -45 41084 -35 43156
rect -2230 41070 -35 41084
rect 35 43156 2230 43170
rect 35 43120 2170 43156
rect 35 41120 85 43120
rect 2085 41120 2170 43120
rect 35 41084 2170 41120
rect 2220 41084 2230 43156
rect 35 41070 2230 41084
rect -2230 40996 -35 41010
rect -2230 40960 -95 40996
rect -2230 38960 -2180 40960
rect -180 38960 -95 40960
rect -2230 38924 -95 38960
rect -45 38924 -35 40996
rect -2230 38910 -35 38924
rect 35 40996 2230 41010
rect 35 40960 2170 40996
rect 35 38960 85 40960
rect 2085 38960 2170 40960
rect 35 38924 2170 38960
rect 2220 38924 2230 40996
rect 35 38910 2230 38924
rect -2230 38836 -35 38850
rect -2230 38800 -95 38836
rect -2230 36800 -2180 38800
rect -180 36800 -95 38800
rect -2230 36764 -95 36800
rect -45 36764 -35 38836
rect -2230 36750 -35 36764
rect 35 38836 2230 38850
rect 35 38800 2170 38836
rect 35 36800 85 38800
rect 2085 36800 2170 38800
rect 35 36764 2170 36800
rect 2220 36764 2230 38836
rect 35 36750 2230 36764
rect -2230 36676 -35 36690
rect -2230 36640 -95 36676
rect -2230 34640 -2180 36640
rect -180 34640 -95 36640
rect -2230 34604 -95 34640
rect -45 34604 -35 36676
rect -2230 34590 -35 34604
rect 35 36676 2230 36690
rect 35 36640 2170 36676
rect 35 34640 85 36640
rect 2085 34640 2170 36640
rect 35 34604 2170 34640
rect 2220 34604 2230 36676
rect 35 34590 2230 34604
rect -2230 34516 -35 34530
rect -2230 34480 -95 34516
rect -2230 32480 -2180 34480
rect -180 32480 -95 34480
rect -2230 32444 -95 32480
rect -45 32444 -35 34516
rect -2230 32430 -35 32444
rect 35 34516 2230 34530
rect 35 34480 2170 34516
rect 35 32480 85 34480
rect 2085 32480 2170 34480
rect 35 32444 2170 32480
rect 2220 32444 2230 34516
rect 35 32430 2230 32444
rect -2230 32356 -35 32370
rect -2230 32320 -95 32356
rect -2230 30320 -2180 32320
rect -180 30320 -95 32320
rect -2230 30284 -95 30320
rect -45 30284 -35 32356
rect -2230 30270 -35 30284
rect 35 32356 2230 32370
rect 35 32320 2170 32356
rect 35 30320 85 32320
rect 2085 30320 2170 32320
rect 35 30284 2170 30320
rect 2220 30284 2230 32356
rect 35 30270 2230 30284
rect -2230 30196 -35 30210
rect -2230 30160 -95 30196
rect -2230 28160 -2180 30160
rect -180 28160 -95 30160
rect -2230 28124 -95 28160
rect -45 28124 -35 30196
rect -2230 28110 -35 28124
rect 35 30196 2230 30210
rect 35 30160 2170 30196
rect 35 28160 85 30160
rect 2085 28160 2170 30160
rect 35 28124 2170 28160
rect 2220 28124 2230 30196
rect 35 28110 2230 28124
rect -2230 28036 -35 28050
rect -2230 28000 -95 28036
rect -2230 26000 -2180 28000
rect -180 26000 -95 28000
rect -2230 25964 -95 26000
rect -45 25964 -35 28036
rect -2230 25950 -35 25964
rect 35 28036 2230 28050
rect 35 28000 2170 28036
rect 35 26000 85 28000
rect 2085 26000 2170 28000
rect 35 25964 2170 26000
rect 2220 25964 2230 28036
rect 35 25950 2230 25964
rect -2230 25876 -35 25890
rect -2230 25840 -95 25876
rect -2230 23840 -2180 25840
rect -180 23840 -95 25840
rect -2230 23804 -95 23840
rect -45 23804 -35 25876
rect -2230 23790 -35 23804
rect 35 25876 2230 25890
rect 35 25840 2170 25876
rect 35 23840 85 25840
rect 2085 23840 2170 25840
rect 35 23804 2170 23840
rect 2220 23804 2230 25876
rect 35 23790 2230 23804
rect -2230 23716 -35 23730
rect -2230 23680 -95 23716
rect -2230 21680 -2180 23680
rect -180 21680 -95 23680
rect -2230 21644 -95 21680
rect -45 21644 -35 23716
rect -2230 21630 -35 21644
rect 35 23716 2230 23730
rect 35 23680 2170 23716
rect 35 21680 85 23680
rect 2085 21680 2170 23680
rect 35 21644 2170 21680
rect 2220 21644 2230 23716
rect 35 21630 2230 21644
rect -2230 21556 -35 21570
rect -2230 21520 -95 21556
rect -2230 19520 -2180 21520
rect -180 19520 -95 21520
rect -2230 19484 -95 19520
rect -45 19484 -35 21556
rect -2230 19470 -35 19484
rect 35 21556 2230 21570
rect 35 21520 2170 21556
rect 35 19520 85 21520
rect 2085 19520 2170 21520
rect 35 19484 2170 19520
rect 2220 19484 2230 21556
rect 35 19470 2230 19484
rect -2230 19396 -35 19410
rect -2230 19360 -95 19396
rect -2230 17360 -2180 19360
rect -180 17360 -95 19360
rect -2230 17324 -95 17360
rect -45 17324 -35 19396
rect -2230 17310 -35 17324
rect 35 19396 2230 19410
rect 35 19360 2170 19396
rect 35 17360 85 19360
rect 2085 17360 2170 19360
rect 35 17324 2170 17360
rect 2220 17324 2230 19396
rect 35 17310 2230 17324
rect -2230 17236 -35 17250
rect -2230 17200 -95 17236
rect -2230 15200 -2180 17200
rect -180 15200 -95 17200
rect -2230 15164 -95 15200
rect -45 15164 -35 17236
rect -2230 15150 -35 15164
rect 35 17236 2230 17250
rect 35 17200 2170 17236
rect 35 15200 85 17200
rect 2085 15200 2170 17200
rect 35 15164 2170 15200
rect 2220 15164 2230 17236
rect 35 15150 2230 15164
rect -2230 15076 -35 15090
rect -2230 15040 -95 15076
rect -2230 13040 -2180 15040
rect -180 13040 -95 15040
rect -2230 13004 -95 13040
rect -45 13004 -35 15076
rect -2230 12990 -35 13004
rect 35 15076 2230 15090
rect 35 15040 2170 15076
rect 35 13040 85 15040
rect 2085 13040 2170 15040
rect 35 13004 2170 13040
rect 2220 13004 2230 15076
rect 35 12990 2230 13004
rect -2230 12916 -35 12930
rect -2230 12880 -95 12916
rect -2230 10880 -2180 12880
rect -180 10880 -95 12880
rect -2230 10844 -95 10880
rect -45 10844 -35 12916
rect -2230 10830 -35 10844
rect 35 12916 2230 12930
rect 35 12880 2170 12916
rect 35 10880 85 12880
rect 2085 10880 2170 12880
rect 35 10844 2170 10880
rect 2220 10844 2230 12916
rect 35 10830 2230 10844
rect -2230 10756 -35 10770
rect -2230 10720 -95 10756
rect -2230 8720 -2180 10720
rect -180 8720 -95 10720
rect -2230 8684 -95 8720
rect -45 8684 -35 10756
rect -2230 8670 -35 8684
rect 35 10756 2230 10770
rect 35 10720 2170 10756
rect 35 8720 85 10720
rect 2085 8720 2170 10720
rect 35 8684 2170 8720
rect 2220 8684 2230 10756
rect 35 8670 2230 8684
rect -2230 8596 -35 8610
rect -2230 8560 -95 8596
rect -2230 6560 -2180 8560
rect -180 6560 -95 8560
rect -2230 6524 -95 6560
rect -45 6524 -35 8596
rect -2230 6510 -35 6524
rect 35 8596 2230 8610
rect 35 8560 2170 8596
rect 35 6560 85 8560
rect 2085 6560 2170 8560
rect 35 6524 2170 6560
rect 2220 6524 2230 8596
rect 35 6510 2230 6524
rect -2230 6436 -35 6450
rect -2230 6400 -95 6436
rect -2230 4400 -2180 6400
rect -180 4400 -95 6400
rect -2230 4364 -95 4400
rect -45 4364 -35 6436
rect -2230 4350 -35 4364
rect 35 6436 2230 6450
rect 35 6400 2170 6436
rect 35 4400 85 6400
rect 2085 4400 2170 6400
rect 35 4364 2170 4400
rect 2220 4364 2230 6436
rect 35 4350 2230 4364
rect -2230 4276 -35 4290
rect -2230 4240 -95 4276
rect -2230 2240 -2180 4240
rect -180 2240 -95 4240
rect -2230 2204 -95 2240
rect -45 2204 -35 4276
rect -2230 2190 -35 2204
rect 35 4276 2230 4290
rect 35 4240 2170 4276
rect 35 2240 85 4240
rect 2085 2240 2170 4240
rect 35 2204 2170 2240
rect 2220 2204 2230 4276
rect 35 2190 2230 2204
rect -2230 2116 -35 2130
rect -2230 2080 -95 2116
rect -2230 80 -2180 2080
rect -180 80 -95 2080
rect -2230 44 -95 80
rect -45 44 -35 2116
rect -2230 30 -35 44
rect 35 2116 2230 2130
rect 35 2080 2170 2116
rect 35 80 85 2080
rect 2085 80 2170 2080
rect 35 44 2170 80
rect 2220 44 2230 2116
rect 35 30 2230 44
rect -2230 -44 -35 -30
rect -2230 -80 -95 -44
rect -2230 -2080 -2180 -80
rect -180 -2080 -95 -80
rect -2230 -2116 -95 -2080
rect -45 -2116 -35 -44
rect -2230 -2130 -35 -2116
rect 35 -44 2230 -30
rect 35 -80 2170 -44
rect 35 -2080 85 -80
rect 2085 -2080 2170 -80
rect 35 -2116 2170 -2080
rect 2220 -2116 2230 -44
rect 35 -2130 2230 -2116
rect -2230 -2204 -35 -2190
rect -2230 -2240 -95 -2204
rect -2230 -4240 -2180 -2240
rect -180 -4240 -95 -2240
rect -2230 -4276 -95 -4240
rect -45 -4276 -35 -2204
rect -2230 -4290 -35 -4276
rect 35 -2204 2230 -2190
rect 35 -2240 2170 -2204
rect 35 -4240 85 -2240
rect 2085 -4240 2170 -2240
rect 35 -4276 2170 -4240
rect 2220 -4276 2230 -2204
rect 35 -4290 2230 -4276
rect -2230 -4364 -35 -4350
rect -2230 -4400 -95 -4364
rect -2230 -6400 -2180 -4400
rect -180 -6400 -95 -4400
rect -2230 -6436 -95 -6400
rect -45 -6436 -35 -4364
rect -2230 -6450 -35 -6436
rect 35 -4364 2230 -4350
rect 35 -4400 2170 -4364
rect 35 -6400 85 -4400
rect 2085 -6400 2170 -4400
rect 35 -6436 2170 -6400
rect 2220 -6436 2230 -4364
rect 35 -6450 2230 -6436
rect -2230 -6524 -35 -6510
rect -2230 -6560 -95 -6524
rect -2230 -8560 -2180 -6560
rect -180 -8560 -95 -6560
rect -2230 -8596 -95 -8560
rect -45 -8596 -35 -6524
rect -2230 -8610 -35 -8596
rect 35 -6524 2230 -6510
rect 35 -6560 2170 -6524
rect 35 -8560 85 -6560
rect 2085 -8560 2170 -6560
rect 35 -8596 2170 -8560
rect 2220 -8596 2230 -6524
rect 35 -8610 2230 -8596
rect -2230 -8684 -35 -8670
rect -2230 -8720 -95 -8684
rect -2230 -10720 -2180 -8720
rect -180 -10720 -95 -8720
rect -2230 -10756 -95 -10720
rect -45 -10756 -35 -8684
rect -2230 -10770 -35 -10756
rect 35 -8684 2230 -8670
rect 35 -8720 2170 -8684
rect 35 -10720 85 -8720
rect 2085 -10720 2170 -8720
rect 35 -10756 2170 -10720
rect 2220 -10756 2230 -8684
rect 35 -10770 2230 -10756
rect -2230 -10844 -35 -10830
rect -2230 -10880 -95 -10844
rect -2230 -12880 -2180 -10880
rect -180 -12880 -95 -10880
rect -2230 -12916 -95 -12880
rect -45 -12916 -35 -10844
rect -2230 -12930 -35 -12916
rect 35 -10844 2230 -10830
rect 35 -10880 2170 -10844
rect 35 -12880 85 -10880
rect 2085 -12880 2170 -10880
rect 35 -12916 2170 -12880
rect 2220 -12916 2230 -10844
rect 35 -12930 2230 -12916
rect -2230 -13004 -35 -12990
rect -2230 -13040 -95 -13004
rect -2230 -15040 -2180 -13040
rect -180 -15040 -95 -13040
rect -2230 -15076 -95 -15040
rect -45 -15076 -35 -13004
rect -2230 -15090 -35 -15076
rect 35 -13004 2230 -12990
rect 35 -13040 2170 -13004
rect 35 -15040 85 -13040
rect 2085 -15040 2170 -13040
rect 35 -15076 2170 -15040
rect 2220 -15076 2230 -13004
rect 35 -15090 2230 -15076
rect -2230 -15164 -35 -15150
rect -2230 -15200 -95 -15164
rect -2230 -17200 -2180 -15200
rect -180 -17200 -95 -15200
rect -2230 -17236 -95 -17200
rect -45 -17236 -35 -15164
rect -2230 -17250 -35 -17236
rect 35 -15164 2230 -15150
rect 35 -15200 2170 -15164
rect 35 -17200 85 -15200
rect 2085 -17200 2170 -15200
rect 35 -17236 2170 -17200
rect 2220 -17236 2230 -15164
rect 35 -17250 2230 -17236
rect -2230 -17324 -35 -17310
rect -2230 -17360 -95 -17324
rect -2230 -19360 -2180 -17360
rect -180 -19360 -95 -17360
rect -2230 -19396 -95 -19360
rect -45 -19396 -35 -17324
rect -2230 -19410 -35 -19396
rect 35 -17324 2230 -17310
rect 35 -17360 2170 -17324
rect 35 -19360 85 -17360
rect 2085 -19360 2170 -17360
rect 35 -19396 2170 -19360
rect 2220 -19396 2230 -17324
rect 35 -19410 2230 -19396
rect -2230 -19484 -35 -19470
rect -2230 -19520 -95 -19484
rect -2230 -21520 -2180 -19520
rect -180 -21520 -95 -19520
rect -2230 -21556 -95 -21520
rect -45 -21556 -35 -19484
rect -2230 -21570 -35 -21556
rect 35 -19484 2230 -19470
rect 35 -19520 2170 -19484
rect 35 -21520 85 -19520
rect 2085 -21520 2170 -19520
rect 35 -21556 2170 -21520
rect 2220 -21556 2230 -19484
rect 35 -21570 2230 -21556
rect -2230 -21644 -35 -21630
rect -2230 -21680 -95 -21644
rect -2230 -23680 -2180 -21680
rect -180 -23680 -95 -21680
rect -2230 -23716 -95 -23680
rect -45 -23716 -35 -21644
rect -2230 -23730 -35 -23716
rect 35 -21644 2230 -21630
rect 35 -21680 2170 -21644
rect 35 -23680 85 -21680
rect 2085 -23680 2170 -21680
rect 35 -23716 2170 -23680
rect 2220 -23716 2230 -21644
rect 35 -23730 2230 -23716
rect -2230 -23804 -35 -23790
rect -2230 -23840 -95 -23804
rect -2230 -25840 -2180 -23840
rect -180 -25840 -95 -23840
rect -2230 -25876 -95 -25840
rect -45 -25876 -35 -23804
rect -2230 -25890 -35 -25876
rect 35 -23804 2230 -23790
rect 35 -23840 2170 -23804
rect 35 -25840 85 -23840
rect 2085 -25840 2170 -23840
rect 35 -25876 2170 -25840
rect 2220 -25876 2230 -23804
rect 35 -25890 2230 -25876
rect -2230 -25964 -35 -25950
rect -2230 -26000 -95 -25964
rect -2230 -28000 -2180 -26000
rect -180 -28000 -95 -26000
rect -2230 -28036 -95 -28000
rect -45 -28036 -35 -25964
rect -2230 -28050 -35 -28036
rect 35 -25964 2230 -25950
rect 35 -26000 2170 -25964
rect 35 -28000 85 -26000
rect 2085 -28000 2170 -26000
rect 35 -28036 2170 -28000
rect 2220 -28036 2230 -25964
rect 35 -28050 2230 -28036
rect -2230 -28124 -35 -28110
rect -2230 -28160 -95 -28124
rect -2230 -30160 -2180 -28160
rect -180 -30160 -95 -28160
rect -2230 -30196 -95 -30160
rect -45 -30196 -35 -28124
rect -2230 -30210 -35 -30196
rect 35 -28124 2230 -28110
rect 35 -28160 2170 -28124
rect 35 -30160 85 -28160
rect 2085 -30160 2170 -28160
rect 35 -30196 2170 -30160
rect 2220 -30196 2230 -28124
rect 35 -30210 2230 -30196
rect -2230 -30284 -35 -30270
rect -2230 -30320 -95 -30284
rect -2230 -32320 -2180 -30320
rect -180 -32320 -95 -30320
rect -2230 -32356 -95 -32320
rect -45 -32356 -35 -30284
rect -2230 -32370 -35 -32356
rect 35 -30284 2230 -30270
rect 35 -30320 2170 -30284
rect 35 -32320 85 -30320
rect 2085 -32320 2170 -30320
rect 35 -32356 2170 -32320
rect 2220 -32356 2230 -30284
rect 35 -32370 2230 -32356
rect -2230 -32444 -35 -32430
rect -2230 -32480 -95 -32444
rect -2230 -34480 -2180 -32480
rect -180 -34480 -95 -32480
rect -2230 -34516 -95 -34480
rect -45 -34516 -35 -32444
rect -2230 -34530 -35 -34516
rect 35 -32444 2230 -32430
rect 35 -32480 2170 -32444
rect 35 -34480 85 -32480
rect 2085 -34480 2170 -32480
rect 35 -34516 2170 -34480
rect 2220 -34516 2230 -32444
rect 35 -34530 2230 -34516
rect -2230 -34604 -35 -34590
rect -2230 -34640 -95 -34604
rect -2230 -36640 -2180 -34640
rect -180 -36640 -95 -34640
rect -2230 -36676 -95 -36640
rect -45 -36676 -35 -34604
rect -2230 -36690 -35 -36676
rect 35 -34604 2230 -34590
rect 35 -34640 2170 -34604
rect 35 -36640 85 -34640
rect 2085 -36640 2170 -34640
rect 35 -36676 2170 -36640
rect 2220 -36676 2230 -34604
rect 35 -36690 2230 -36676
rect -2230 -36764 -35 -36750
rect -2230 -36800 -95 -36764
rect -2230 -38800 -2180 -36800
rect -180 -38800 -95 -36800
rect -2230 -38836 -95 -38800
rect -45 -38836 -35 -36764
rect -2230 -38850 -35 -38836
rect 35 -36764 2230 -36750
rect 35 -36800 2170 -36764
rect 35 -38800 85 -36800
rect 2085 -38800 2170 -36800
rect 35 -38836 2170 -38800
rect 2220 -38836 2230 -36764
rect 35 -38850 2230 -38836
rect -2230 -38924 -35 -38910
rect -2230 -38960 -95 -38924
rect -2230 -40960 -2180 -38960
rect -180 -40960 -95 -38960
rect -2230 -40996 -95 -40960
rect -45 -40996 -35 -38924
rect -2230 -41010 -35 -40996
rect 35 -38924 2230 -38910
rect 35 -38960 2170 -38924
rect 35 -40960 85 -38960
rect 2085 -40960 2170 -38960
rect 35 -40996 2170 -40960
rect 2220 -40996 2230 -38924
rect 35 -41010 2230 -40996
rect -2230 -41084 -35 -41070
rect -2230 -41120 -95 -41084
rect -2230 -43120 -2180 -41120
rect -180 -43120 -95 -41120
rect -2230 -43156 -95 -43120
rect -45 -43156 -35 -41084
rect -2230 -43170 -35 -43156
rect 35 -41084 2230 -41070
rect 35 -41120 2170 -41084
rect 35 -43120 85 -41120
rect 2085 -43120 2170 -41120
rect 35 -43156 2170 -43120
rect 2220 -43156 2230 -41084
rect 35 -43170 2230 -43156
rect -2230 -43244 -35 -43230
rect -2230 -43280 -95 -43244
rect -2230 -45280 -2180 -43280
rect -180 -45280 -95 -43280
rect -2230 -45316 -95 -45280
rect -45 -45316 -35 -43244
rect -2230 -45330 -35 -45316
rect 35 -43244 2230 -43230
rect 35 -43280 2170 -43244
rect 35 -45280 85 -43280
rect 2085 -45280 2170 -43280
rect 35 -45316 2170 -45280
rect 2220 -45316 2230 -43244
rect 35 -45330 2230 -45316
rect -2230 -45404 -35 -45390
rect -2230 -45440 -95 -45404
rect -2230 -47440 -2180 -45440
rect -180 -47440 -95 -45440
rect -2230 -47476 -95 -47440
rect -45 -47476 -35 -45404
rect -2230 -47490 -35 -47476
rect 35 -45404 2230 -45390
rect 35 -45440 2170 -45404
rect 35 -47440 85 -45440
rect 2085 -47440 2170 -45440
rect 35 -47476 2170 -47440
rect 2220 -47476 2230 -45404
rect 35 -47490 2230 -47476
rect -2230 -47564 -35 -47550
rect -2230 -47600 -95 -47564
rect -2230 -49600 -2180 -47600
rect -180 -49600 -95 -47600
rect -2230 -49636 -95 -49600
rect -45 -49636 -35 -47564
rect -2230 -49650 -35 -49636
rect 35 -47564 2230 -47550
rect 35 -47600 2170 -47564
rect 35 -49600 85 -47600
rect 2085 -49600 2170 -47600
rect 35 -49636 2170 -49600
rect 2220 -49636 2230 -47564
rect 35 -49650 2230 -49636
rect -2230 -49724 -35 -49710
rect -2230 -49760 -95 -49724
rect -2230 -51760 -2180 -49760
rect -180 -51760 -95 -49760
rect -2230 -51796 -95 -51760
rect -45 -51796 -35 -49724
rect -2230 -51810 -35 -51796
rect 35 -49724 2230 -49710
rect 35 -49760 2170 -49724
rect 35 -51760 85 -49760
rect 2085 -51760 2170 -49760
rect 35 -51796 2170 -51760
rect 2220 -51796 2230 -49724
rect 35 -51810 2230 -51796
rect -2230 -51884 -35 -51870
rect -2230 -51920 -95 -51884
rect -2230 -53920 -2180 -51920
rect -180 -53920 -95 -51920
rect -2230 -53956 -95 -53920
rect -45 -53956 -35 -51884
rect -2230 -53970 -35 -53956
rect 35 -51884 2230 -51870
rect 35 -51920 2170 -51884
rect 35 -53920 85 -51920
rect 2085 -53920 2170 -51920
rect 35 -53956 2170 -53920
rect 2220 -53956 2230 -51884
rect 35 -53970 2230 -53956
rect -2230 -54044 -35 -54030
rect -2230 -54080 -95 -54044
rect -2230 -56080 -2180 -54080
rect -180 -56080 -95 -54080
rect -2230 -56116 -95 -56080
rect -45 -56116 -35 -54044
rect -2230 -56130 -35 -56116
rect 35 -54044 2230 -54030
rect 35 -54080 2170 -54044
rect 35 -56080 85 -54080
rect 2085 -56080 2170 -54080
rect 35 -56116 2170 -56080
rect 2220 -56116 2230 -54044
rect 35 -56130 2230 -56116
rect -2230 -56204 -35 -56190
rect -2230 -56240 -95 -56204
rect -2230 -58240 -2180 -56240
rect -180 -58240 -95 -56240
rect -2230 -58276 -95 -58240
rect -45 -58276 -35 -56204
rect -2230 -58290 -35 -58276
rect 35 -56204 2230 -56190
rect 35 -56240 2170 -56204
rect 35 -58240 85 -56240
rect 2085 -58240 2170 -56240
rect 35 -58276 2170 -58240
rect 2220 -58276 2230 -56204
rect 35 -58290 2230 -58276
rect -2230 -58364 -35 -58350
rect -2230 -58400 -95 -58364
rect -2230 -60400 -2180 -58400
rect -180 -60400 -95 -58400
rect -2230 -60436 -95 -60400
rect -45 -60436 -35 -58364
rect -2230 -60450 -35 -60436
rect 35 -58364 2230 -58350
rect 35 -58400 2170 -58364
rect 35 -60400 85 -58400
rect 2085 -60400 2170 -58400
rect 35 -60436 2170 -60400
rect 2220 -60436 2230 -58364
rect 35 -60450 2230 -60436
<< viatp >>
rect -95 58364 -45 60436
rect 2170 58364 2220 60436
rect -95 56204 -45 58276
rect 2170 56204 2220 58276
rect -95 54044 -45 56116
rect 2170 54044 2220 56116
rect -95 51884 -45 53956
rect 2170 51884 2220 53956
rect -95 49724 -45 51796
rect 2170 49724 2220 51796
rect -95 47564 -45 49636
rect 2170 47564 2220 49636
rect -95 45404 -45 47476
rect 2170 45404 2220 47476
rect -95 43244 -45 45316
rect 2170 43244 2220 45316
rect -95 41084 -45 43156
rect 2170 41084 2220 43156
rect -95 38924 -45 40996
rect 2170 38924 2220 40996
rect -95 36764 -45 38836
rect 2170 36764 2220 38836
rect -95 34604 -45 36676
rect 2170 34604 2220 36676
rect -95 32444 -45 34516
rect 2170 32444 2220 34516
rect -95 30284 -45 32356
rect 2170 30284 2220 32356
rect -95 28124 -45 30196
rect 2170 28124 2220 30196
rect -95 25964 -45 28036
rect 2170 25964 2220 28036
rect -95 23804 -45 25876
rect 2170 23804 2220 25876
rect -95 21644 -45 23716
rect 2170 21644 2220 23716
rect -95 19484 -45 21556
rect 2170 19484 2220 21556
rect -95 17324 -45 19396
rect 2170 17324 2220 19396
rect -95 15164 -45 17236
rect 2170 15164 2220 17236
rect -95 13004 -45 15076
rect 2170 13004 2220 15076
rect -95 10844 -45 12916
rect 2170 10844 2220 12916
rect -95 8684 -45 10756
rect 2170 8684 2220 10756
rect -95 6524 -45 8596
rect 2170 6524 2220 8596
rect -95 4364 -45 6436
rect 2170 4364 2220 6436
rect -95 2204 -45 4276
rect 2170 2204 2220 4276
rect -95 44 -45 2116
rect 2170 44 2220 2116
rect -95 -2116 -45 -44
rect 2170 -2116 2220 -44
rect -95 -4276 -45 -2204
rect 2170 -4276 2220 -2204
rect -95 -6436 -45 -4364
rect 2170 -6436 2220 -4364
rect -95 -8596 -45 -6524
rect 2170 -8596 2220 -6524
rect -95 -10756 -45 -8684
rect 2170 -10756 2220 -8684
rect -95 -12916 -45 -10844
rect 2170 -12916 2220 -10844
rect -95 -15076 -45 -13004
rect 2170 -15076 2220 -13004
rect -95 -17236 -45 -15164
rect 2170 -17236 2220 -15164
rect -95 -19396 -45 -17324
rect 2170 -19396 2220 -17324
rect -95 -21556 -45 -19484
rect 2170 -21556 2220 -19484
rect -95 -23716 -45 -21644
rect 2170 -23716 2220 -21644
rect -95 -25876 -45 -23804
rect 2170 -25876 2220 -23804
rect -95 -28036 -45 -25964
rect 2170 -28036 2220 -25964
rect -95 -30196 -45 -28124
rect 2170 -30196 2220 -28124
rect -95 -32356 -45 -30284
rect 2170 -32356 2220 -30284
rect -95 -34516 -45 -32444
rect 2170 -34516 2220 -32444
rect -95 -36676 -45 -34604
rect 2170 -36676 2220 -34604
rect -95 -38836 -45 -36764
rect 2170 -38836 2220 -36764
rect -95 -40996 -45 -38924
rect 2170 -40996 2220 -38924
rect -95 -43156 -45 -41084
rect 2170 -43156 2220 -41084
rect -95 -45316 -45 -43244
rect 2170 -45316 2220 -43244
rect -95 -47476 -45 -45404
rect 2170 -47476 2220 -45404
rect -95 -49636 -45 -47564
rect 2170 -49636 2220 -47564
rect -95 -51796 -45 -49724
rect 2170 -51796 2220 -49724
rect -95 -53956 -45 -51884
rect 2170 -53956 2220 -51884
rect -95 -56116 -45 -54044
rect 2170 -56116 2220 -54044
rect -95 -58276 -45 -56204
rect 2170 -58276 2220 -56204
rect -95 -60436 -45 -58364
rect 2170 -60436 2220 -58364
<< metaltp >>
rect -1215 60385 -1145 60480
rect -105 60436 -35 60480
rect -1215 58225 -1145 58415
rect -105 58364 -95 60436
rect -45 58364 -35 60436
rect 1050 60385 1120 60480
rect 2160 60436 2230 60480
rect -105 58276 -35 58364
rect -1215 56065 -1145 56255
rect -105 56204 -95 58276
rect -45 56204 -35 58276
rect 1050 58225 1120 58415
rect 2160 58364 2170 60436
rect 2220 58364 2230 60436
rect 2160 58276 2230 58364
rect -105 56116 -35 56204
rect -1215 53905 -1145 54095
rect -105 54044 -95 56116
rect -45 54044 -35 56116
rect 1050 56065 1120 56255
rect 2160 56204 2170 58276
rect 2220 56204 2230 58276
rect 2160 56116 2230 56204
rect -105 53956 -35 54044
rect -1215 51745 -1145 51935
rect -105 51884 -95 53956
rect -45 51884 -35 53956
rect 1050 53905 1120 54095
rect 2160 54044 2170 56116
rect 2220 54044 2230 56116
rect 2160 53956 2230 54044
rect -105 51796 -35 51884
rect -1215 49585 -1145 49775
rect -105 49724 -95 51796
rect -45 49724 -35 51796
rect 1050 51745 1120 51935
rect 2160 51884 2170 53956
rect 2220 51884 2230 53956
rect 2160 51796 2230 51884
rect -105 49636 -35 49724
rect -1215 47425 -1145 47615
rect -105 47564 -95 49636
rect -45 47564 -35 49636
rect 1050 49585 1120 49775
rect 2160 49724 2170 51796
rect 2220 49724 2230 51796
rect 2160 49636 2230 49724
rect -105 47476 -35 47564
rect -1215 45265 -1145 45455
rect -105 45404 -95 47476
rect -45 45404 -35 47476
rect 1050 47425 1120 47615
rect 2160 47564 2170 49636
rect 2220 47564 2230 49636
rect 2160 47476 2230 47564
rect -105 45316 -35 45404
rect -1215 43105 -1145 43295
rect -105 43244 -95 45316
rect -45 43244 -35 45316
rect 1050 45265 1120 45455
rect 2160 45404 2170 47476
rect 2220 45404 2230 47476
rect 2160 45316 2230 45404
rect -105 43156 -35 43244
rect -1215 40945 -1145 41135
rect -105 41084 -95 43156
rect -45 41084 -35 43156
rect 1050 43105 1120 43295
rect 2160 43244 2170 45316
rect 2220 43244 2230 45316
rect 2160 43156 2230 43244
rect -105 40996 -35 41084
rect -1215 38785 -1145 38975
rect -105 38924 -95 40996
rect -45 38924 -35 40996
rect 1050 40945 1120 41135
rect 2160 41084 2170 43156
rect 2220 41084 2230 43156
rect 2160 40996 2230 41084
rect -105 38836 -35 38924
rect -1215 36625 -1145 36815
rect -105 36764 -95 38836
rect -45 36764 -35 38836
rect 1050 38785 1120 38975
rect 2160 38924 2170 40996
rect 2220 38924 2230 40996
rect 2160 38836 2230 38924
rect -105 36676 -35 36764
rect -1215 34465 -1145 34655
rect -105 34604 -95 36676
rect -45 34604 -35 36676
rect 1050 36625 1120 36815
rect 2160 36764 2170 38836
rect 2220 36764 2230 38836
rect 2160 36676 2230 36764
rect -105 34516 -35 34604
rect -1215 32305 -1145 32495
rect -105 32444 -95 34516
rect -45 32444 -35 34516
rect 1050 34465 1120 34655
rect 2160 34604 2170 36676
rect 2220 34604 2230 36676
rect 2160 34516 2230 34604
rect -105 32356 -35 32444
rect -1215 30145 -1145 30335
rect -105 30284 -95 32356
rect -45 30284 -35 32356
rect 1050 32305 1120 32495
rect 2160 32444 2170 34516
rect 2220 32444 2230 34516
rect 2160 32356 2230 32444
rect -105 30196 -35 30284
rect -1215 27985 -1145 28175
rect -105 28124 -95 30196
rect -45 28124 -35 30196
rect 1050 30145 1120 30335
rect 2160 30284 2170 32356
rect 2220 30284 2230 32356
rect 2160 30196 2230 30284
rect -105 28036 -35 28124
rect -1215 25825 -1145 26015
rect -105 25964 -95 28036
rect -45 25964 -35 28036
rect 1050 27985 1120 28175
rect 2160 28124 2170 30196
rect 2220 28124 2230 30196
rect 2160 28036 2230 28124
rect -105 25876 -35 25964
rect -1215 23665 -1145 23855
rect -105 23804 -95 25876
rect -45 23804 -35 25876
rect 1050 25825 1120 26015
rect 2160 25964 2170 28036
rect 2220 25964 2230 28036
rect 2160 25876 2230 25964
rect -105 23716 -35 23804
rect -1215 21505 -1145 21695
rect -105 21644 -95 23716
rect -45 21644 -35 23716
rect 1050 23665 1120 23855
rect 2160 23804 2170 25876
rect 2220 23804 2230 25876
rect 2160 23716 2230 23804
rect -105 21556 -35 21644
rect -1215 19345 -1145 19535
rect -105 19484 -95 21556
rect -45 19484 -35 21556
rect 1050 21505 1120 21695
rect 2160 21644 2170 23716
rect 2220 21644 2230 23716
rect 2160 21556 2230 21644
rect -105 19396 -35 19484
rect -1215 17185 -1145 17375
rect -105 17324 -95 19396
rect -45 17324 -35 19396
rect 1050 19345 1120 19535
rect 2160 19484 2170 21556
rect 2220 19484 2230 21556
rect 2160 19396 2230 19484
rect -105 17236 -35 17324
rect -1215 15025 -1145 15215
rect -105 15164 -95 17236
rect -45 15164 -35 17236
rect 1050 17185 1120 17375
rect 2160 17324 2170 19396
rect 2220 17324 2230 19396
rect 2160 17236 2230 17324
rect -105 15076 -35 15164
rect -1215 12865 -1145 13055
rect -105 13004 -95 15076
rect -45 13004 -35 15076
rect 1050 15025 1120 15215
rect 2160 15164 2170 17236
rect 2220 15164 2230 17236
rect 2160 15076 2230 15164
rect -105 12916 -35 13004
rect -1215 10705 -1145 10895
rect -105 10844 -95 12916
rect -45 10844 -35 12916
rect 1050 12865 1120 13055
rect 2160 13004 2170 15076
rect 2220 13004 2230 15076
rect 2160 12916 2230 13004
rect -105 10756 -35 10844
rect -1215 8545 -1145 8735
rect -105 8684 -95 10756
rect -45 8684 -35 10756
rect 1050 10705 1120 10895
rect 2160 10844 2170 12916
rect 2220 10844 2230 12916
rect 2160 10756 2230 10844
rect -105 8596 -35 8684
rect -1215 6385 -1145 6575
rect -105 6524 -95 8596
rect -45 6524 -35 8596
rect 1050 8545 1120 8735
rect 2160 8684 2170 10756
rect 2220 8684 2230 10756
rect 2160 8596 2230 8684
rect -105 6436 -35 6524
rect -1215 4225 -1145 4415
rect -105 4364 -95 6436
rect -45 4364 -35 6436
rect 1050 6385 1120 6575
rect 2160 6524 2170 8596
rect 2220 6524 2230 8596
rect 2160 6436 2230 6524
rect -105 4276 -35 4364
rect -1215 2065 -1145 2255
rect -105 2204 -95 4276
rect -45 2204 -35 4276
rect 1050 4225 1120 4415
rect 2160 4364 2170 6436
rect 2220 4364 2230 6436
rect 2160 4276 2230 4364
rect -105 2116 -35 2204
rect -1215 -95 -1145 95
rect -105 44 -95 2116
rect -45 44 -35 2116
rect 1050 2065 1120 2255
rect 2160 2204 2170 4276
rect 2220 2204 2230 4276
rect 2160 2116 2230 2204
rect -105 -44 -35 44
rect -1215 -2255 -1145 -2065
rect -105 -2116 -95 -44
rect -45 -2116 -35 -44
rect 1050 -95 1120 95
rect 2160 44 2170 2116
rect 2220 44 2230 2116
rect 2160 -44 2230 44
rect -105 -2204 -35 -2116
rect -1215 -4415 -1145 -4225
rect -105 -4276 -95 -2204
rect -45 -4276 -35 -2204
rect 1050 -2255 1120 -2065
rect 2160 -2116 2170 -44
rect 2220 -2116 2230 -44
rect 2160 -2204 2230 -2116
rect -105 -4364 -35 -4276
rect -1215 -6575 -1145 -6385
rect -105 -6436 -95 -4364
rect -45 -6436 -35 -4364
rect 1050 -4415 1120 -4225
rect 2160 -4276 2170 -2204
rect 2220 -4276 2230 -2204
rect 2160 -4364 2230 -4276
rect -105 -6524 -35 -6436
rect -1215 -8735 -1145 -8545
rect -105 -8596 -95 -6524
rect -45 -8596 -35 -6524
rect 1050 -6575 1120 -6385
rect 2160 -6436 2170 -4364
rect 2220 -6436 2230 -4364
rect 2160 -6524 2230 -6436
rect -105 -8684 -35 -8596
rect -1215 -10895 -1145 -10705
rect -105 -10756 -95 -8684
rect -45 -10756 -35 -8684
rect 1050 -8735 1120 -8545
rect 2160 -8596 2170 -6524
rect 2220 -8596 2230 -6524
rect 2160 -8684 2230 -8596
rect -105 -10844 -35 -10756
rect -1215 -13055 -1145 -12865
rect -105 -12916 -95 -10844
rect -45 -12916 -35 -10844
rect 1050 -10895 1120 -10705
rect 2160 -10756 2170 -8684
rect 2220 -10756 2230 -8684
rect 2160 -10844 2230 -10756
rect -105 -13004 -35 -12916
rect -1215 -15215 -1145 -15025
rect -105 -15076 -95 -13004
rect -45 -15076 -35 -13004
rect 1050 -13055 1120 -12865
rect 2160 -12916 2170 -10844
rect 2220 -12916 2230 -10844
rect 2160 -13004 2230 -12916
rect -105 -15164 -35 -15076
rect -1215 -17375 -1145 -17185
rect -105 -17236 -95 -15164
rect -45 -17236 -35 -15164
rect 1050 -15215 1120 -15025
rect 2160 -15076 2170 -13004
rect 2220 -15076 2230 -13004
rect 2160 -15164 2230 -15076
rect -105 -17324 -35 -17236
rect -1215 -19535 -1145 -19345
rect -105 -19396 -95 -17324
rect -45 -19396 -35 -17324
rect 1050 -17375 1120 -17185
rect 2160 -17236 2170 -15164
rect 2220 -17236 2230 -15164
rect 2160 -17324 2230 -17236
rect -105 -19484 -35 -19396
rect -1215 -21695 -1145 -21505
rect -105 -21556 -95 -19484
rect -45 -21556 -35 -19484
rect 1050 -19535 1120 -19345
rect 2160 -19396 2170 -17324
rect 2220 -19396 2230 -17324
rect 2160 -19484 2230 -19396
rect -105 -21644 -35 -21556
rect -1215 -23855 -1145 -23665
rect -105 -23716 -95 -21644
rect -45 -23716 -35 -21644
rect 1050 -21695 1120 -21505
rect 2160 -21556 2170 -19484
rect 2220 -21556 2230 -19484
rect 2160 -21644 2230 -21556
rect -105 -23804 -35 -23716
rect -1215 -26015 -1145 -25825
rect -105 -25876 -95 -23804
rect -45 -25876 -35 -23804
rect 1050 -23855 1120 -23665
rect 2160 -23716 2170 -21644
rect 2220 -23716 2230 -21644
rect 2160 -23804 2230 -23716
rect -105 -25964 -35 -25876
rect -1215 -28175 -1145 -27985
rect -105 -28036 -95 -25964
rect -45 -28036 -35 -25964
rect 1050 -26015 1120 -25825
rect 2160 -25876 2170 -23804
rect 2220 -25876 2230 -23804
rect 2160 -25964 2230 -25876
rect -105 -28124 -35 -28036
rect -1215 -30335 -1145 -30145
rect -105 -30196 -95 -28124
rect -45 -30196 -35 -28124
rect 1050 -28175 1120 -27985
rect 2160 -28036 2170 -25964
rect 2220 -28036 2230 -25964
rect 2160 -28124 2230 -28036
rect -105 -30284 -35 -30196
rect -1215 -32495 -1145 -32305
rect -105 -32356 -95 -30284
rect -45 -32356 -35 -30284
rect 1050 -30335 1120 -30145
rect 2160 -30196 2170 -28124
rect 2220 -30196 2230 -28124
rect 2160 -30284 2230 -30196
rect -105 -32444 -35 -32356
rect -1215 -34655 -1145 -34465
rect -105 -34516 -95 -32444
rect -45 -34516 -35 -32444
rect 1050 -32495 1120 -32305
rect 2160 -32356 2170 -30284
rect 2220 -32356 2230 -30284
rect 2160 -32444 2230 -32356
rect -105 -34604 -35 -34516
rect -1215 -36815 -1145 -36625
rect -105 -36676 -95 -34604
rect -45 -36676 -35 -34604
rect 1050 -34655 1120 -34465
rect 2160 -34516 2170 -32444
rect 2220 -34516 2230 -32444
rect 2160 -34604 2230 -34516
rect -105 -36764 -35 -36676
rect -1215 -38975 -1145 -38785
rect -105 -38836 -95 -36764
rect -45 -38836 -35 -36764
rect 1050 -36815 1120 -36625
rect 2160 -36676 2170 -34604
rect 2220 -36676 2230 -34604
rect 2160 -36764 2230 -36676
rect -105 -38924 -35 -38836
rect -1215 -41135 -1145 -40945
rect -105 -40996 -95 -38924
rect -45 -40996 -35 -38924
rect 1050 -38975 1120 -38785
rect 2160 -38836 2170 -36764
rect 2220 -38836 2230 -36764
rect 2160 -38924 2230 -38836
rect -105 -41084 -35 -40996
rect -1215 -43295 -1145 -43105
rect -105 -43156 -95 -41084
rect -45 -43156 -35 -41084
rect 1050 -41135 1120 -40945
rect 2160 -40996 2170 -38924
rect 2220 -40996 2230 -38924
rect 2160 -41084 2230 -40996
rect -105 -43244 -35 -43156
rect -1215 -45455 -1145 -45265
rect -105 -45316 -95 -43244
rect -45 -45316 -35 -43244
rect 1050 -43295 1120 -43105
rect 2160 -43156 2170 -41084
rect 2220 -43156 2230 -41084
rect 2160 -43244 2230 -43156
rect -105 -45404 -35 -45316
rect -1215 -47615 -1145 -47425
rect -105 -47476 -95 -45404
rect -45 -47476 -35 -45404
rect 1050 -45455 1120 -45265
rect 2160 -45316 2170 -43244
rect 2220 -45316 2230 -43244
rect 2160 -45404 2230 -45316
rect -105 -47564 -35 -47476
rect -1215 -49775 -1145 -49585
rect -105 -49636 -95 -47564
rect -45 -49636 -35 -47564
rect 1050 -47615 1120 -47425
rect 2160 -47476 2170 -45404
rect 2220 -47476 2230 -45404
rect 2160 -47564 2230 -47476
rect -105 -49724 -35 -49636
rect -1215 -51935 -1145 -51745
rect -105 -51796 -95 -49724
rect -45 -51796 -35 -49724
rect 1050 -49775 1120 -49585
rect 2160 -49636 2170 -47564
rect 2220 -49636 2230 -47564
rect 2160 -49724 2230 -49636
rect -105 -51884 -35 -51796
rect -1215 -54095 -1145 -53905
rect -105 -53956 -95 -51884
rect -45 -53956 -35 -51884
rect 1050 -51935 1120 -51745
rect 2160 -51796 2170 -49724
rect 2220 -51796 2230 -49724
rect 2160 -51884 2230 -51796
rect -105 -54044 -35 -53956
rect -1215 -56255 -1145 -56065
rect -105 -56116 -95 -54044
rect -45 -56116 -35 -54044
rect 1050 -54095 1120 -53905
rect 2160 -53956 2170 -51884
rect 2220 -53956 2230 -51884
rect 2160 -54044 2230 -53956
rect -105 -56204 -35 -56116
rect -1215 -58415 -1145 -58225
rect -105 -58276 -95 -56204
rect -45 -58276 -35 -56204
rect 1050 -56255 1120 -56065
rect 2160 -56116 2170 -54044
rect 2220 -56116 2230 -54044
rect 2160 -56204 2230 -56116
rect -105 -58364 -35 -58276
rect -1215 -60480 -1145 -60385
rect -105 -60436 -95 -58364
rect -45 -60436 -35 -58364
rect 1050 -58415 1120 -58225
rect 2160 -58276 2170 -56204
rect 2220 -58276 2230 -56204
rect 2160 -58364 2230 -58276
rect -105 -60480 -35 -60436
rect 1050 -60480 1120 -60385
rect 2160 -60436 2170 -58364
rect 2220 -60436 2230 -58364
rect 2160 -60480 2230 -60436
<< properties >>
string parameters w 20.00 l 20.00 val 413.6 carea 1.00 cperi 0.17 nx 2 ny 56 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string gencell cmm5t
string library efxh018
<< end >>
